MZP      ��  �       @                                     � �	�!�L�!��This program must be run under Win32
$7                                                                                                                                                                                                                                                                                                                                                                                                        PE  L �dM        � #                         @                      0	                                                    	                                                                                                         .text                                `.data                             @  �.rsrc     	     	                @  @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �ZW>          @  �   `  �   �  �
   � �    �     �    �ZW>          8 �   P �    �ZW>       y  h �y  � �y  � �    �ZW>      d    � �   � �   � �   � �	    �
   ( �   @ �   X �   p �   � �   � �   � �   � �   � �     �    �   0 �   H �   ` �   x �   � �   � �   � �   � �    � �!    �&     �'   8 �B   P �E   h �F   � �G   � �H   � �I   � �J   � �R   � �S   	 �T   (	 �U   @	 �X   X	 �Y   p	 �\   �	 �]   �	 �^   �	 �_   �	 �e   �	 �f    
 �g   
 �h   0
 �i   H
 �j   `
 �k   x
 �l   �
 �m   �
 �n   �
 �o   �
 �p   �
 �q    �r     �s   8 �t   P �w   h �x   � �~   � �   � ��   � ��   � ��   � ��    ��   ( ��   @ �  X �  p �  � �  � �  � �  � �  � �    ��   ��  0 ��  H ��  ` ��  x ��  � ��  � ��  � ��  � ��  � ��   ��    ��  8 ��  P ��  h ��  � ��  � ��  � ��  � ��  � �   � �    �ZW>    (   0 � �> �( �X �@ �| �X �� �p �� �� �� �� �� �� �, �� �N �� �| �  �� � �� �0 �� �H � �` �: �x �Z �� �� �� �� �� �� �� � �� �* � �Z �  �l �8 �� �P �� �h �� �� �� �� �  �� �8  �� �\  �� ��  �� ��  � ��  �( ��  �@ �! �X �,! �p �J! �� ��! �� ��! �� �    �ZW>       y  � �    �ZW>          � �    �ZW>                �ZW>               �ZW>                �ZW>         0      �ZW>         @      �ZW>         P      �ZW>         `      �ZW>         p      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>                �ZW>               �ZW>                �ZW>         0      �ZW>         @      �ZW>         P      �ZW>         `      �ZW>         p      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>                �ZW>               �ZW>                �ZW>         0      �ZW>         @      �ZW>         P      �ZW>         `      �ZW>         p      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>                �ZW>               �ZW>                �ZW>         0      �ZW>         @      �ZW>         P      �ZW>         `      �ZW>         p      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>                �ZW>               �ZW>                �ZW>         0      �ZW>         @      �ZW>         P      �ZW>         `      �ZW>         p      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>                �ZW>               �ZW>                �ZW>         0      �ZW>         @      �ZW>         P      �ZW>         `      �ZW>         p      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>         �      �ZW>                �ZW>               �ZW>                �ZW>         0      �ZW>         @      �ZW>         P      �ZW>         `      �ZW>         p      �ZW>         �      �ZW>           �      �ZW>           �      �ZW>           �      �ZW>           �      �ZW>           �      �ZW>           �      �ZW>           �      �ZW>                  �ZW>                 �ZW>                  �ZW>           0      �ZW>           @      �ZW>           P      �ZW>           `      �ZW>           p      �ZW>           �      �ZW>           �      �ZW>           �      �ZW>           �      �ZW>           �      �ZW>           �      �ZW>           �      �ZW>           �      �ZW>                  �ZW>                 �ZW>                  �ZW>           0      �ZW>           @      �ZW>           P      �ZW>           `      �ZW>           p      �ZW>           �      �ZW>           �      �ZW>           �      �ZW>           �      �ZW>           �      �ZW>           �      �ZW>           �      �ZW>           �      �ZW>                  �ZW>               �ZW>            �1  4          3  �           �3  �           |4  l          �5  D          ,7  �          �V  �=          L�  J          ��  b          ��            �  v          ��            ��  ^          �  D          L�  �          �  (          <�  6          t�  �          ��  ^          T�  ~          ��  �          ��  �          ��  �          H�  |          ��  �          ��  x          ��  B          @�  �          4�  �          ��  J          H  |           �  �          � �          X �          D �            `          x |          �$ &          3           ,; &          T<           \C �          H �          �\ 0           e �          �f �          \h .          �i �          <p           L} ,          x �          4� R          �� n          �� v           p� *          �� �          T� �          ,� �          ̌ �          �� �          @� �          �� �          ė           ܙ v          T� "          x� 8           �� �           �� �          0�           D� N          �� X          � h          T� (          |� l           � �           �� x           ,� >           l� J          �� �          D� �          � �          ļ �           p� �          4� d          �� �          T�           X� �           4� x          �� ,          �� �          �� B          � �          �� 8          �� �           �� �           0� �          �� p          X� �          4� �          �� j          ,� �          �� X           �           ,� *          X�           \�            l� �         �� �          � �          �� �          �� .
          �� �          �� *          �            �          � �
          T( �           + /          0? bf          ��           �� 6
          � �          �� �          p� �          $� �          �  T          < L(          �+ �          T4 �
          ? ��          � ��          D� �          � �           x I          l� `          ̚ �          P� T          �� �>          �� �|          �a R          �� �          ��           �� �S          �	 �          0$	 �          �)	 "           �)	 D           D V C L A L  T A B O U T D I A L O G  T A U T H E N T I C A T E F O R M  T C L E A N U P D I A L O G  T C O N S O L E D I A L O G  T C O P Y D I A L O G  T C O P Y P A R A M C U S T O M D I A L O G  T C O P Y P A R A M P R E S E T D I A L O G  T C O P Y P A R A M S F R A M E  T C R E A T E D I R E C T O R Y D I A L O G  T C U S T O M C O M M A N D D I A L O G  T C U S T O M D I A L O G  T C U S T O M S C P E X P L O R E R F O R M  T E D I T O R F O R M  T E D I T O R P R E F E R E N C E S D I A L O G  T F I L E F I N D D I A L O G  T F I L E S Y S T E M I N F O D I A L O G  T F U L L S Y N C H R O N I Z E D I A L O G  T G E N E R A L S E T T I N G S F R A M E  T I M P O R T S E S S I O N S D I A L O G  T L I C E N S E D I A L O G  T L O C A T I O N P R O F I L E S D I A L O G  T L O G F O R M  T L O G G I N G F R A M E  T L O G I N D I A L O G  T N O N V I S U A L D A T A M O D U L E  T O P E N D I R E C T O R Y D I A L O G  T P R E F E R E N C E S D I A L O G  T P R O G R E S S F O R M  T P R O P E R T I E S D I A L O G  T R E M O T E T R A N S F E R D I A L O G  T R I G H T S E X T F R A M E  T R I G H T S F R A M E  T S C P C O M M A N D E R F O R M  T S C P E X P L O R E R F O R M  T S E L E C T M A S K D I A L O G  T S Y M L I N K D I A L O G  T S Y N C H R O N I Z E C H E C K L I S T D I A L O G  T S Y N C H R O N I Z E D I A L O G  T S Y N C H R O N I Z E P R O G R E S S F O R M     (       @                                ���                                  8   0   p   `   �   �  �  �  �  �  �  �  �  �  �                                 ����������������������������������������������������?��?��?� �?�  ?�  �p ���������������������������  (                �                       ��� �  �  ��  �H  �x  �H  ��  �d  ��  �)  �9  �  ��  �|  �   �   �  �  x  0�  �  �         !              �  �  ?�  (      
         P                         �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ��� �����  �����  �www�  �  �  ����  �  �  �����  �����  �����          (   '                                    �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                     ����� ����  ����� ����� ������ ����� ���� ����� ����� ������ ����� ���� ����� ����� ������ ����� ���� ����� ����� ������ ����� ���� ����� ����� ������ ����� ����  �����                     (   !            �                         �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ��� �����������������   ������������wwww�   ������������w�ww�   ������� ���x�ww�   �������  ������w�   ������� ���x�w�   ��������� ���w���   ��������� ��wwx��   ������������www��   ������������wwww�   �����������������     US e r v e r n s   v � r d n y c k e l   h i t t a d e s   i n t e   i   c a c h e n .   D e t   f i n n s   i n g e n   g a r a n t i   a t t   s e r v e r n   � r   d e n   d u   t r o r   d e t   � r . 
 
 S e r v e r n s   % s   f i n g e r a v t r y c k s n y c k e l   � r : 
 % s 
 
 O m   d u   l i t a r   p �   v � r d e n ,   t r y c k   J a .   F � r   a t t   a n s l u t a   u t a n   a t t   l � g g a   t i l l   v � r d n y c k e l   i   c a c h e n ,   t r y c k   N e j .   F � r   a t t   � v e r g e   a n s l u t n i n g e n   t r y c k   A v b r y t . 
 
 F o r t s � t t   a n s l u t a   o c h   l � g g a   t i l l   v � r d n y c k e l   i   c a c h e n ? �V A R N I N G   -   E V E N T U E L L T   S � K E R H E T S H � L ! 
 
 S e r v e r n s   v � r d n y c k e l   s t � m m e r   i n t e   m e d   d e n   s o m   W i n S C P   h a r   i   c a c h e n .   D e t   b e t y d e r   a t t   a n t i n g e n   s e r v e r n s   a d m i n i s t r a t � r   h a r   b y t t   v � r d n y c k e l ,   s e r v e r n   f � r i n s t � l l e r   o l i k a   n y c k e l   u n d e r   v i s s a   o m s t � n d i g h e t e r ,   e l l e r   a t t   d u   f a k t i s k t   h a r   a n s l u t i t   t i l l   e n   d a t o r   s o m   l � t s a s   v a r a   s e r v e r n . 
 
 D e n   n y a   % s   f i n g e r a v t r y c k s n y c k e l n   � r : 
 % s 
 
 O m   d u   f � r v � n t a d e   d e n n a   � n d r i n g ,   l i t a   p �   d e n   n y a   n y c k e l   o c h   v i l l   f o r t s � t t a   a n s l u t a ,   a n t i n g e n   t r y c k   U p p d a t e r a   f � r   a t t   u p p d a t e r a   c a c h e ,   e l l e r   t r y c k   L � g g   t i l l   f � r   a t t   l � g g a   t i l l   d e n   n y a   n y c k e l   t i l l   c a c h e n   m e d a n   d e   g a m l a   b e h � l l s .   O m   d u   v i l l   f o r t s � t t a   a n s l u t a   m e n   u t a n   u p p d a t e r a   c a c h e n ,   t r y c k   H o p p a   � v e r .   O m   d u   v i l l   � v e r g e   a n s l u t n i n g   t o t a l t ,   t r y c k   A v b r y t .   T r y c k a   A v b r y t   � r   d e t   E N D A   g a r a n t e r a t   s � k r a   v a l e t . 
 0D u   l a d d a r   e n   S S H - 2   p r i v a t   n y c k e l   s o m   h a r   e t t   g a m m a l t   f i l f o r m a t .   D e t   i n n e b � r   a t t   d i n   n y c k e l f i l   i n t e   � r   h e l t   s � k e r   f � r   m a n i p u l e r i n g s f � r s � k .   V i   r e k o m m e n d e r a r   d i g   a t t   k o n v e r t e r a   d i n   n y c k e l   t i l l   d e t   n y a   f o r m a t e t . 
 
 D u   k a n   u t f � r a   d e n   h � r   k o n v e r t e r i n g e n   g e n o m   a t t   l a d d a   f i l e n   i   P u T T Y g e n   o c h   s e d a n   s p a r a   d e n   i g e n . � H e l p   [   < k o m m a n d o >   [   < k o m m a n d o 2 >   . . .   ] 
     V i s a r   l i s t a   p �   k o m m a n d o n   o m   i n g a   p a r a m e t e r a r   a n g e s . 
     V i s a r   h j � l p   o m   e t t   k o m m a n d o   o m   d e t   a n g e s . 
 a l i a s : 
     m a n 
 e x e m p e l : 
     h e l p 
     h e l p   l s 
 D e x i t 
     S t � n g e r   a l l a   s e s s i o n e r   o c h   a v s l u t a r   p r o g r a m m e t . 
 a l i a s : 
     b y e 
 To p e n   < s t o r e d   s e s s i o n > 
 o p e n   [   s f t p | s c p | f t p : / /   ] [   < u s e r >   [   : p a s s w o r d   ]   @   ]   < h o s t >   [   : < p o r t >   ] 
     U p p r � t t a r   a n s l u t n i n g   t i l l   g i v e n   v � r d .   A n v � n d   a n t i n g e n   n a m n e t   p �   d e n   l a g r a d e 
     s e s s i o n e n   e l l e r   a n g e   v � r d ,   a n v � n d a r n a m n ,   p o r t   o c h   p r o t o k o l l   d i r e k t . 
 s w i t c h e s : 
     - p r i v a t e k e y = < k e y >     P r i v a t e   n y c k e l f i l 
     - t i m e o u t = < s e c >           S e r v e r s v a r   t i m e o u t 
     - h o s t k e y = < f i n g e r p r i n t >   F i n g e r a v t r y c k   f � r   s e r v e r n s   v � r d n y c k e l   ( e n d a s t   S F T P   o c h   S C P ) . 
     - c e r t i f i c a t e = < f i n g e r p r i n t >   F i n g e r a v t r y c k   f � r   S S L / T L S   c e r t i f i k a t   ( e n d a s t   F T P S ) 
     - p a s s i v e                       P a s s i v t   l � g e   ( e n d a s t   F T P   p r o t o k o l l ) 
     - i m p l i c i t                     I m p l i c i t   T L S / S S L   ( e n d a s t   F T P S   p r o t o k o l l ) 
     - e x p l i c i t s s l               E x p l i c i t   S S L   ( e n d a s t   F T P S   p r o t o k o l l ) 
     - e x p l i c i t t l s               E x p l i c i t   T L S   ( e n d a s t   F T P S   p r o t o k o l l ) 
 e x a m p l e s : 
     o p e n 
     o p e n   s f t p : / / m a r t i n @ e x a m p l e . c o m : 2 2 2 2   - p r i v a t e k e y = m y k e y . p p k 
     o p e n   m a r t i n @ e x a m p l e . c o m 
     o p e n   e x a m p l e . c o m 
 � c l o s e   [   < s e s s i o n >   ] 
     S t � n g e r   s e s s i o n   s p e c i f i c e r a d   m e d   s i t t   n u m m e r .   O m   s e s s i o n s n u m r e t   i n t e   � r 
     s p e c i f i c e r a d ,   s t � n g s   d e n   a k t u e l l a   s e s s i o n e n . 
 e x e m p e l : 
     c l o s e 
     c l o s e   1 
 � s e s s i o n   [   < s e s s i o n >   ] 
     G � r   s e s s i o n e n   s p e c i f i c e r a d   m e d   e t t   n u m m e r   a k t i v .   O m   e t t   s e s s i o n s n u m m e r 
     i n t e   � r   s p e c i f i c e r a d ,   l i s t a s   a n s l u t n a   s e s s i o n e r . 
 e x e m p e l : 
     s e s s i o n 
     s e s s i o n   1 
 ; p w d 
     V i s a r   a k t u e l l   f j � r r k a t a l o g   f � r   d e n   a k t i v a   s e s s i o n e n . 
 � c d   [   < k a t a l o g >   ] 
     � n d r a r   a k t u e l l   k a t a l o g   p �   s e r v e r n   i   d e n   a k t i v a   s e s s i o n e n . 
     O m   e n   k a t a l o g   i n t e   a n g e s ,   a n v � n d s   h e m k a t a l o g e n . 
 e x e m p e l : 
     c d   / h o m e / m a r t i n 
     c d 
 l s   [   < k a t a l o g >   ] / [   < j o k e r t e c k e n > ] 
     V i s a r   i n n e h � l l e t   i   a n g i v e n   f j � r r k a t a l o g .   O m   k a t a l o g   
   i n t e   a n g e s ,   v i s a s   i n n e h � l l e t   i   a k t u e l l   k a t a l o g . 
     N � r   j o k e r t e c k e n   h a r   a n g e t t s ,   t o l k a s   d e t   s o m   e n   g r u p p   f i l e r   s k a   l i s t a s . 
   A n n a r s   l i s t a s   a l l a   f i l e r . 
 a s l i a s : 
     d i r 
 e x e m p e l : 
     l s 
     l s   / h o m e / m a r t i n 
 @ l p w d 
     V i s a r   a k t u e l l   l o k a l   k a t a l o g   ( g � l l e r   f � r   a l l a   s e s s i o n e r ) . 
 J l c d   < k a t a l o g > 
     B y t e r   l o k a l   k a t a l o g   f � r   a l l a   s e s s i o n e r . 
 e x e m p e l : 
     c d   d : \ 
 l l s   [   < k a t a l o g >   ] \ [   < j o k e r t e c k e n >   ] 
     V i s a r   i n n e h � l l e t   i   a n g i v e n   l o k a l   k a t a l o g .   O m   k a t a l o g   
     i n t e   a n g e s ,   v i s a s   i n n e h � l l e t   i   a k t u e l l   k a t a l o g . 
     N � r   j o k e r t e c k e n   h a r   a n g e t t s ,   t o l k a s   d e t   s o m   e n   g r u p p   f i l e r   s k a   l i s t a s . 
   A n n a r s   l i s t a s   a l l a   f i l e r . 
 e x e m p e l : 
     l l s 
     l l s   d : \ 
 r m   < f i l >   [   < f i l 2 >   . . .   ] 
     R a d e r a r   e n   e l l e r   f l e r a   f j � r r f i l e r .   O m   f j � r r p a p p e r s k o r g e n   � r 
     k o n f i g u r e r a d ,   f l y t t a s   f i l e n   d i t   i s t � l l e t   f � r   a t t   r a d e r a s . 
     F i l n a m n   k a n   e r s � t t a s   a v   j o k e r t e c k e n   f � r   a t t   v � l j a   f l e r a   f i l e r . 
 e x e m p e l : 
     r m   i n d e x . h t m l 
     r m   i n d e x . h t m l   a b o u t . h t m l 
     r m   * . h t m l 
 � r m d i r   < k a t a l o g >   [   < k a t a l o g 2 >   . . .   ] 
     R a d e r a r   e n   e l l e r   f l e r a   f j � r r k a t a l o g e r .   O m   f j � r r p a p p e r s k o r g e n   � r 
   k o n f i g u r e r a d ,   f l y t t a s   k a t a l o g e n   d i t   i s t � l l e t   f � r   a t t   r a d e r a s . 
 e x e m p e l : 
     r m d i r   p u b l i c _ h t m l 
  m v   < f i l >   [   < f i l 2 >   . . .   ]   [   < k a t a l o g > /   ] [   < n y t t n a m n >   ] 
     F l y t t a r   e l l e r   b y t e r   n a m n   p �   e n   e l l e r   f l e r a   f j � r r f i l e r .   M � l k a t a l o g e n   e l l e r   n y t t 
     n a m n   e l l e r   b � d a   m � s t e   a n g e s .   M � l k a t a l o g e n   m � s t e   a v s l u t a s   m e d   
     s n e d s t r e c k .   O p e r a t i o n s m a s k   k a n   a n v � n d a s   i s t � l l e t   f � r   n y t t   n a m n . 
     F i l n a m n   k a n   b y t a s   u t   m o t   j o k e r t e c k e n   f � r   a t t   v � l j a   f l e r a   f i l e r . 
 a l i a s : 
     r e n a m e 
 e x e m p e l : 
     m v   i n d e x . h t m l   p u b l c _ h t m l / 
     m v   i n d e x . h t m l   a b o u t . * 
     m v   i n d e x . h t m l   p u b l i c _ h t m l / a b o u t . * 
     m v   p u b l i c _ h t m l / i n d e x . h t m l   p u b l i c _ h t m l / a b o u t . h t m l   / h o m e / m a r t i n / * . b a k 
     m v   * . h t m l   / h o m e / b a c k u p / * . b a k 
 :c h m o d   < m e t o d >   < f i l >   [   < f i l 2 >   . . .   ] 
     � n d r a r   r � t t i g h e t e r n a   p �   e n   e l l e r   f l e r a   f j � r r f i l e r .   M e t o d   k a n   a n g e s 
     s o m   t r e -   e l l e r   f y r s i f f r i g a   o k t a l a   n u m m e r . 
     F i l n a m n   k a n   b y t a s   u t   m o t   j o k e r t e c k e n   f � r   a t t   v � l j a   f l e r a   f i l e r . 
 e x e m p e l : 
     c h m o d   6 4 4   i n d e x . h t m l   a b o u t . h t m l 
     c h m o d   1 7 0 0   / h o m e / m a r t i n / p u b l i c _ h t m l 
     c h m o d   6 4 4   * . h t m l 
 m l n   < m � l >   < s y m l � n k > 
     S k a p a r   s y m b o l i s k   f j � r r l � n k . 
 a l i a s : 
     s y m l i n k 
 e x e m p e l : 
     l n   / h o m e / m a r t i n / p u b l i c _ h t m l   w w w 
 D m k d i r   < k a t a l o g > 
     S k a p a r   f j � r r k a t a l o g . 
 e x e m p e l : 
     m k d i r   p u b l i c _ h t m l 
 :g e t   < f i l >   [   [   < f i l 2 >   . . .   ]   < k a t a l o g > \ [   < n y t t _ n a m n >   ]   ] 
     L a d d a r   n e r   e n   e l l e r   f l e r   f i l e r   f r � n   f j � r r k a t a l o g   t i l l   l o k a l   k a t a l o g . 
     O m   e n d a s t   e n   p a r a m e t e r   � r   a n g i v e n   l a d d a s   f i l e n   t i l l   e n   l o k a l   a r b e t s k a t a l o g . 
     O m   f l e r a   p a r a m e t r a r   a n g e s ,   a n g e r   a l l a 
   f � r u t o m   d e n   s i s t a   v i l k e n   g r u p p   f i l e r   s o m   s k a   l a d d a s   n e r .   D e n   s i s t a   p a r a m e t e r n   a n g e r   m � l e t 
   p �   l o k a l   k a t a l o g   o c h   e v e n t u e l l   o p e r a t i o n s m a s k   f � r   a t t   l a g r a   f i l ( e r )   u n d e r 
     a n n a t   n a m n .   M � l k a t a l o g e n   m � s t e   s l u t a   m e d   e t t   o m v � n t   s n e d s t r e c k . 
     F i l n a m n   k a n   e r s � t t a s   m e d   j o k e r t e c k e n   f � r   a t t   m a r k e r a   f l e r a   f i l e r . 
     F � r   a t t   l a d d a   n e r   f l e r   f i l e r   t i l l   a k t u e l l   a r b e t s k a t a l o g   a n v � n d   ' . \ '   s o m   d e n   
   s i s t a   p a r a m e t e r n . 
     A n v � n d   ' o p t i o n '   k o m m a n d o t   f � r   a t t   s t � l l a   i n   � v e r f � r i n g s a l t e r n a t i v . 
 a l i a s : 
     r e c v 
 s w i t c h e s : 
     - d e l e t e                   R a d e r a r   k � l l a   f � r   f j � r r f i l ( e r )   e f t e r   � v e r f � r i n g   
     - r e s u m e                   � t e r u p p t a   � v e r f � r i n g   o m   m � j l i g t   ( S F T P   o c h   F T P   p r o t o k o l l e n   e n d a s t ) 
     - a p p e n d                   B i f o g a   f i l   t i l l   s l u t e t   a v   m � l f i l   ( S F T P   p r o t o k o l l   e n d a s t ) 
     - p r e s e r v e t i m e       B e v a r a   t i d s s t � m p e l 
     - n o p r e s e r v e t i m e   B e v a r a   i n t e   t i d s s t � m p e l 
     - s p e e d = < k i b p s >     B e g r � n s a   � v e r f � r i n g s h a s t i g h e t 
 e f f e c t i v e   o p t i o n s : 
     t r a n s f e r ,   c o n f i r m ,   e x c l u d e ,   i n c l u d e ,   r e c o n n e c t t i m e 
 e x a m p l e s : 
     g e t   i n d e x . h t m l 
     g e t   - d e l e t e   i n d e x . h t m l   a b o u t . h t m l   . \ 
     g e t   i n d e x . h t m l   a b o u t . h t m l   d : \ w w w \ 
     g e t   p u b l i c _ h t m l / i n d e x . h t m l   d : \ w w w \ a b o u t . * 
     g e t   * . h t m l   * . p n g   d : \ w w w \ * . b a k 
 �p u t   < f i l >   [   [   < f i l 2 >   . . .   ]   < k a t a l o g > / [   < n y t t _ n a m n >   ]   ] 
     L a d d a r   u p p   e n   e l l e r   f l e r a   f i l e r   f r � n   l o k a l   k a t a l o g   t i l l   f j � r r k a t a l o g . 
     O m   e n d a s t   e n   p a r a m e t e r   a n g e s   l a d d a s   f i l e n   t i l l   e n 
   f j � r r a r b e t s k a t a l o g .   O m   f l e r   p a r a m e t r a r   a n g e s ,   a n g e   a l l a   f � r u t o m   d e n   s i s t a 
     v i l k e n   g r u p p   f i l e r   s o m   s k a   l a d d a s   u p p .   D e n   s i s t a   p a r a m e t e r n   a n g e r   m � l e t 
     p �   f j � r r k a t a l o g   o c h   e v e n t u e l l   o p e r a t i o n s m a s k   f � r   a t t   l a g r a   f i l ( e r )   u n d e r 
     a n n a t   n a m n .   M � l k a t a l o g e n   m � s t e   s l u t a   m e d   e t t   s n e d s t r e c k .   
     F i l n a m n   k a n   e r s � t t a s   m e d   j o k e r t e c k e n   f � r   a t t   m a r k e r a   f l e r a   f i l e r . 
     F � r   a t t   l a d d a   u p p   f l e r a   f i l e r   t i l l   a k t u e l l   a r b e t s k a t a l o g ,   a n v � n d   ' . / '   s o m   d e n 
     s i s t a   p a r a m e t e r n . 
     A n v � n d   ' o p t i o n '   k o m m a n d o t   f � r   a t t   s t � l l a   i n   � v e r f � r i n g s a l t e r n a t i v . 
 a l i a s : 
     s e n d 
 s w i t c h e s : 
     - d e l e t e                           R a d e r a r   k � l l a   f � r   l o k a l   f i l ( e r )   e f t e r   � v e r f � r i n g 
     - r e s u m e                           � t e r u p p t a r   � v e r f � r i n g   o m   m � j l i g t   ( S F T P   o c h   F T P   p r o k o l l e n   e n d a s t ) 
     - a p p e n d                           B i f o g a   f i l   t i l l   s l u t e t   a v   m � l f i l   ( F T P   p r o t o k o l l   e n d a s t ) 
     - p r e s e r v e t i m e               B e v a r a   t i d s s t � m p e l 
     - n o p r e s e r v e t i m e           B e v a r a   i n t e   t i d s s t � m p e l 
     - p e r m i s s i o n s = < m o d e >   A n g e   r � t t i g h e t e r 
     - n o p e r m i s s i o n s             B e v a r a   s t a n d a r d r � t t i g h e t e r 
     - s p e e d = < k i b p s >             B e g r � n s a   � v e r f � r i n g s h a s t i g h e t 
 e f f e c t i v e   o p t i o n s : 
     t r a n s f e r ,   c o n f i r m ,   e x c l u d e ,   i n c l u d e ,   r e c o n n e c t t i m e 
 e x a m p l e s : 
     p u t   i n d e x . h t m l 
     p u t   - d e l e t e   i n d e x . h t m l   a b o u t . h t m l   . / 
     p u t   - p e r m i s s i o n s = 6 4 4   i n d e x . h t m l   a b o u t . h t m l   / h o m e / m a r t i n / p u b l i c _ h t m l / 
     p u t   d : \ w w w \ i n d e x . h t m l   a b o u t . * 
     p u t   * . h t m l   * . p n g   / h o m e / m a r t i n / b a c k u p / * . b a k 
  o p t i o n   [   < a l t e r n a t i v >   [   < v � r d e >   ]   ] 
     O m   i n g a   p a r a m e t r a r   a n g e s ,   v i s a s   a l l a   s c r i p t   a l t e r n a t i v   o c h 
   d e r a s   v � r d e n .   O m   e n d a s t   e n   p a r a m e t e r   a n g e s ,   v i s a s   v � r d e t   f � r   a l t e r n a t i v e t . 
     O m   t v �   p a r a m e t r a r   a n g e s   s � t t   v � r d e t   p �   a l t e r n a t i v e t . 
     U r s p r u n g l i g a   v � r d e n   a v   v i s s a   a l t e r n a t i v   � r   h � m t a d e   f r � n   a p p l i k a t i o n e n s   k o n f i g u r a t i o n , 
     m o d i f i k a t i o n   a v   d e s s a   � n d r a d   d o c k   i n t e   a p p l i k a t i o n e n s 
   k o n f i g u r a t i o n . 
 o p t i o n s   a r e : 
     e c h o           o n | o f f 
                       V � x l a r   e k o   a v   k o m m a n d o   s o m   e x e k v e r a s . 
                       C o m m a n d s   a f f e c t e d :   a l l 
     b a t c h         o n | o f f | a b o r t | c o n t i n u e 
                       V � x l a r   b a t c h   l � g e   ( a l l a   u p p m a n i n g a r   b e s v a r a s   a u t o m a t i s k t 
                       n e g a t i v t ) .   N � r   ' o n ' ,   r e k o m m e n d e r a s   a t t   s � t t a   ' c o n f i r m ' 
                       t i l l   ' o f f '   f � r   a t t   t i l l � t a   � v e r s k r i v n i n g a r .   M e d   ' a b o r t ' ,   s c r i p t   a v b r y t s 
                       n � r   e t t   f e l   i n t r � f f a r .   M e d   ' c o n t i n u e ' ,   a l l a   f e l   i g n o r e r a s . 
                       C o m m a n d s   a f f e c t e d :   n e a r l y   a l l 
     c o n f i r m     o n | o f f 
                       V � x l a r   b e k r � f t e l s e r   ( � v e r s k r i v n i n g ,   e t c . ) . 
                       C o m m a n d s   a f f e c t e d :   g e t ,   p u t 
     t r a n s f e r   b i n a r y | a s c i i | a u t o m a t i c 
                       � v e r f � r i n g s l � g e :   b i n a r y ,   a s c i i   ( t e x t ) ,   a u t o m a t i c   ( b y   e x t e n s i o n ) . 
                       C o m m a n d s   a f f e c t e d :   g e t ,   p u t ,   s y n c h r o n i z e ,   k e e p u p t o d a t e 
     e x c l u d e     c l e a r   |   < m a s k >   [   ;   < m a s k 2 >   . . .   ] 
     i n c l u d e     c l e a r   |   < m a s k >   [   ;   < m a s k 2 >   . . .   ] 
                       S t � l l e r   i n   e x k l u d e r i n g s -   e l l e r   i n k l u d e r i n g s m a s k e r   ( e n d a s t   e n   k a n   v a r a   a k t i v ) . 
                       K a t a l o g e r   p � v e r k a s   o c k s �   ( * /   m a t c h a r   a l l a   k a t a l o g e r ) . 
                       C o m m a n d s   a f f e c t e d :   g e t ,   p u t ,   s y n c h r o n i z e ,   k e e p u p t o d a t e 
     r e c o n n e c t t i m e   o f f   |   < s e c > 
                       T i d s b e g r � n s n i n g   i   s e k u n d e r   f � r   � t e r a n s l u t n i n g   a v   b r u t e n   s e s s i o n . 
                       C o m m a n d s   a f f e c t e d :   g e t ,   p u t ,   s y n c h r o n i z e ,   k e e p u p t o d a t e 
 a l i a s e s : 
     a s c i i   =     o p t i o n   t r a n s f e r   a s c i i 
     b i n a r y   =   o p t i o n   t r a n s f e r   b i n a r y 
 e x a m p l e s : 
     o p t i o n 
     o p t i o n   t r a n s f e r 
     o p t i o n   c o n f i r m   o f f 
     o p t i o n   i n c l u d e   " * . h t m l ;   * / " 
 -s y n c h r o n i z e   l o c a l | r e m o t e | b o t h   [   < l o k a l   k a t a l o g >   [   < f j � r r k a t a l o g >   ]   ] 
     N � r   d e n   f � r s t a   p a r a m e t e r n   � r   ' l o c a l '   s y n k r o n i s e r a s   l o k a l   k a t a l o g   m e d 
   f j � r r k a t a l o g .   N � r   d e n   f � r s t a   p a r a m e t e r n   � r   ' r e m o t e '   s y n k r o n i s e r a s   f j � r r k a t a l o g 
   m e d   l o k a l   k a t a l o g .   N � r   f � r s t a   p a r a m e t e r n   � r   ' b o t h '   s y n k r o n i s e r a s 
   k a t a l o g e r n a   e n   m o t   d e n   a n d r a . 
     N � r   i n g e n   k a t a l o g   a n g e s ,   s y n k r o n i s e r a s   a k t u e l l   a r b e t s k a t a l o g .   
     N o t e r a :   � v e r s k r i v n i n g s b e k r � f t e l s e r   � r   a l l t i d   a v s t � n g d a   f � r   k o m m a n d o t . 
 s w i t c h e s : 
     - d e l e t e                             R a d e r a   f � r � l d r a d e   f i l e r 
     - m i r r o r                             M i r r o r   l � g e   ( s y n k r o n i s e r a s   o c k s �   � l d r e   f i l e r ) . 
                                               I g n o r e r a   f � r   ' b o t h ' . 
     - c r i t e r i a = < c r i t e r i a >   J � m f � r e l s e   k r i t e r i e r .   M � j l i g a   v � r d e n   � r   ' n o n e ' ,   ' t i m e ' , 
                                               ' s i z e '   o c h   ' b o t h ' .   I g n o r e r a s   f � r   ' b o t h '   l � g e . 
     - p e r m i s s i o n s = < m o d e >     A n g e   r � t t i g h e t e r 
     - n o p e r m i s s i o n s               B e v a r a   s t a n d a r d r � t t i g h e t e r 
     - s p e e d = < k i b p s >               B e g r � n s a   � v e r f � r i n g s h a s t i g h e t 
 e f f e c t i v e   o p t i o n s : 
     t r a n s f e r ,   e x c l u d e ,   i n c l u d e ,   r e c o n n e c t t i m e 
 e x a m p l e s : 
     s y n c h r o n i z e   r e m o t e   - d e l e t e 
     s y n c h r o n i z e   b o t h   d : \ w w w   / h o m e / m a r t i n / p u b l i c _ h t m l 
 uk e e p u p t o d a t e   [   < l o k a l   k a t a l o g >   [   < f j � r r k a t a l o g >   ]   ] 
     B e v a k a r   � n d r i n g a r   i   l o k a l   k a t a l o g   o c h   � t e r s p e g l a r   d e   p �   f j � r r k a t a l o g . 
     O m   k a t l o g e r   i n t e   a n g e s ,   a k t u e l l   k a t a l o g   s y n k r o n i s e r a s . 
     F � r   a t t   s l u t a   � v e r v a k n i n g   a v   � n d r i n g a r   t r y c k   C T R L - C . 
     N o t e r a :   M e d d e l a n d e n   o m   � v e r s k r i v n i n g   � r   a l l t i d   a v s t � n g d a   f � r   k o m m a n d o t . 
 s w i t c h e s : 
     - d e l e t e                           R a d e r a   g a m l a   f i l e r 
     - p e r m i s s i o n s = < m o d e >   S � t t   r � t t i g h e t e r 
     - n o p e r m i s s i o n s             B e h � l l   s t a n d a r d r � t t i g h e t e r 
     - s p e e d = < k i b p s >             B e g r � n s a   � v e r f � r i n g s h a s t i g h e t 
 e f f e c t i v e   o p t i o n s : 
     t r a n s f e r ,   e x c l u d e ,   i n c l u d e 
 e x a m p l e s : 
     k e e p u p t o d a t e   - d e l e t e 
     k e e p u p t o d a t e   d : \ w w w   / h o m e / m a r t i n / p u b l i c _ h t m l 
 Wc a l l   < K o m m a n d o > 
     M e d   S F T P   o c h   S C P   p r o t o k o l l e n ,   k � r s   g o d t y c k l i g t   f j � r r s k a l s k o m m a n d o . 
     O m   a k t u e l l   s e s s i o n   i n t e   t i l l � t e r   k � r n i n g   a v   g o d t y c k l i g   f j � r r k o m m a n d o 
     s k i l d a   s k a l s e s s i o n e r   k o m m e r   a t t   � p p n a s   a u t o m a t i s k t . 
     O m   F T P   p r o t o k o l l ,   k � r   e t t   p r o t o k o l l k o m m a n d o . 
     K o m m a n d o t   k a n   i n t e   k r � v a   a n v � n d a r i n p u t . 
 a l i a s : 
     ! 
 e x e m p e l : 
     c a l l   t o u c h   i n d e x . h t m l 
                   
 C O R E _ E R R O R " V � r d n y c k e l n   k u n d e   i n t e   v e r i f i e r a s !  A n s l u t n i n g   m i s s l y c k a d e s .  A v s l u t a d   a v   a n v � n d a r e n .  T a p p a d   a n s l u t n i n g . # K a n   i n t e   h i t t a   k o m m a n d o t s   r e t u r k o d . C K o m m a n d o t   ' % s ' 
 m i s s l y c k a d e s   m e d   r e t u r k o d e n   % d   o c h   f e l m e d d e l a n d e 
 % s . ) K o m m a n d o t   m i s s l y c k a d e s   m e d   r e t u r k o d e n   % d . 7 K o m m a n d o t   ' % s '   m i s s l y c k a d e s   m e d   o g i l t i g   u t m a t n i n g   ' % s ' . = F e l   u p p s t o d   n � r   n a m n e t   p �   a k t u e l l   f j � r r k a t a l o g   s k u l l e   h � m t a s . | F e l   u p p s t o d   n � r   s t a r t m e d d e l a n d e   h o p p a d e s   � v e r .   D i t t   s k a l   � r   a n t a g l i g e n   i n k o m p a t i b e l t   m e d   a p p l i k a t i o n e n   ( B A S H   r e k o m m e n d e r a s ) . ) F e l   u p p s t o d   n � r   k a t a l o g   b y t t e s   t i l l   ' % s ' .     ) F e l   u p p s t o d   n � r   l i s t n i n g   a v   k a t a l o g   ' % s ' . % O v � n t a d   k a t a l o g l i s t n i n g   v i d   r a d   ' % s ' . # F e l a k t i g   r � t t i g h e t s b e s k r i v n i n g   ' % s ' ; F e l   u p p s t o d   n � r   d e n   a l l m � n n a   k o n f i g u r a t i o n e n   s k u l l e   r e n s a s . + F e l   u p p s t o d   n � r   l a g r a d e   s e s s i o n e r   r e n s a d e s . / F e l   u p p s t o d   n � r   f i l   m e d   s l u m p t a l s f r � n   r e n s a d e s . - F e l   u p p s t o d   n � r   c a c h a d e   v � r d n y c k l a r   r e n s a d e s . Q F e l   u p p s t o d   n � r   v a r i a b e l   i n n e h � l l a n d e   r e t u r k o d   a v   s e n a s t e   k o m m a n d o   s k u l l e   h i t t a s . 0 F e l   u p p s t o d   n � r   a n v � n d a r g r u p p e r   s k u l l e   s l � s   u p p .  F i l   e l l e r   m a p p   ' % s '   f i n n s   i n t e . ) K a n   i n t e   h i t t a   a t t r i b u t e n   f � r   f i l e n   ' % s ' .  K a n   i n t e   � p p n a   f i l e n   ' % s ' . ( F e l   u p p s t o d   n � r   f i l e n   ' % s '   s k u l l e   l � s a s . 3 A l l v a r l i g t   f e l   u p p s t o d   v i d   k o p i e r i n g   a v   f i l e n   ' % s ' . 0 F i l k o p i e r i n g e n   t i l l   f j � r r k a t a l o g e n   m i s s l y c k a d e s .   0 F i l k o p i e r i n g e n   f r � n   f j � r r k a t a l o g e n   m i s s l y c k a d e s . % S C P   p r o t o k o l l f e l :   O v � n t a d   r a d b r y t n i n g & S C P   p r o t o k o l l f e l :   F e l a k t i g t   t i d s f o r m a t 2 S C P   p r o t o k o l l f e l :   F e l a k t i g   c o n t r o l   r e c o r d   ( % s ;   % s ) # K o p i e r i n g   a v   f i l   ' % s '   m i s s l y c k a d e s . 1 S C P   p r o t o k o l l f e l :   F e l a k t i g t   f i l b e s k r i v n i n g s f o r m a t  ' % s '   � r   i n g e n   m a p p ! % F e l   u p p s t o d   n � r   m a p p e n   ' % s '   s k a p a d e s .  K a n   i n t e   s k a p a   f i l e n   ' % s ' . * F e l   u p p s t o d   v i d   s k r i v n i n g   t i l l   f i l e n   ' % s ' . * K a n   i n t e   s � t t a   a t t r i b u t e n   t i l l   f i l e n   ' % s ' . + F e l m e d d e l a n d e   m o t t a g e t   f r � n   f j � r r s i d a :   ' % s ' " F e l   v i d   b o r t t a g n i n g   a v   f i l e n   ' % s ' . 7 F e l   u p p s t o d   v i d   l o g g n i n g   o c h   d e n   h a r   d � r f � r   s t � n g t s   a v .  K a n   i n t e   � p p n a   l o g g f i l e n   ' % s ' . 0 F e l   u p p s t o d   n � r   f i l e n   ' % s '   b y t t e   n a m n   t i l l   ' % s ' .     F i l e n   m e d   n a m n   ' % s '   f i n n s   r e d a n . $ K a t a l o g e n   m e d   n a m n   ' % s '   f i n n s   r e d a n . 2 F e l   u p p s t o d   v i d   b y t e   a v   k a t a l o g   t i l l   h e m k a t a l o g e n . ' F e l   u p p s t o d   v i d   r e n s n i n g   a v   a l l a   a l i a s .   ; F e l   u p p s t o d   n � r   n a t i o n e l l a   a n v � n d a r v a r i a b l e r   s k u l l e   r e n s a s . ! O v � n t a d   i n d a t a   f r � n   s e r v e r n :   ' % s ' ( F e l   u p p s t o d   n � r   I N I - f i l e n   s k u l l e   r e n s a s .   6 A u t e n t i s e r i n g s l o g g   ( s e   s e s s i o n s l o g g   f � r   d e t a l j e r ) : 
 % s 
  A u t e n t i s e r i n g   m i s s l y c k a d e s . # A n s l u t n i n g e n   h a r   o v � n t a t   a v s l u t a t s . 1 F e l   u p p s t o d   n � r   n y c k e l n   s p a r a d e s   t i l l   f i l e n   ' % s ' .   ) S e r v e r n   s k i c k a d e   k o m m a n d o t   s l u t s t a t u s   % d . < S F T P   p r o t o k o l l v a r n i n g :   F e l a k t i g   m e d d e l a n d e t y p   v i d   s v a r   ( % d ) .   I S F T P - s e r v e r n s   v e r s i o n   ( % d )   s t � d s   i n t e .   V e r s i o n e r   s o m   s t � d s   � r   % d   t i l l   % d . E S F T P   p r o t o k o l l v a r n i n g :   F e l a k t i g t   m e d d e l a n d e n u m m e r   % d   ( f � r v � n t a d e   % d ) .  O v � n t a d   O K   r e s p o n s .  O v � n t a d   E O F   r e s p o n s . ! F i l e n   e l l e r   k a t a l o g e n   f i n n s   i n t e .  � t k o m s t   n e k a d . . A l l m � n t   f e l   ( s e r v e r n   b o r d e   g e   f e l b e s k r i v n i n g ) . J D � l i g t   m e d d e l a n d e   ( D � l i g t   f o r m a t e r a t   p a k e t   e l l e r   i n k o m p a t i b e l t   p r o t o k o l l ) .  I n g e n   a n s l u t n i n g .  F � r l o r a d   a n s l u t n i n g .   S e r v e r n   s t � d e r   i n t e   o p e r a t i o n e n . = % s 
 F e l k o d :   % d 
 F e l m e d d e l a n d e   f r � n   s e r v e r n % s :   % s 
 B e g � r d   k o d :   % d  O k � n d   s t a t u s k o d . ' F e l   v i d   l � s n i n g   a v   s y m b o l i s k   l � n k   ' % s ' . 4 S e r v e r n   r e t u r n e r a d e   t o m   l i s t n i n g   f � r   k a t a l o g e n   ' % s ' . 6 M o t t o g   S S H _ F X P _ N A M E   p a k e t   m e d   n o l l   e l l e r   f l e r a   p o s t e r .   + K a n   i n t e   f �   d e n   v e r k l i g a   s � k v � g e n   f � r   ' % s ' . ) K a n   i n t e   � n d r a   e g e n s k a p e r   f � r   f i l e n   ' % s ' . F K a n   i n t e   i n i t i a l i s e r a   S F T P - p r o t o k o l l e t .   K � r   v � r d d a t o r n   e n   S F T P - s e r v e r ? " K a n   i n t e   l � s a   t i d s z o n s i n f o r m a t i o n .  K a n   i n t e   s k a p a   f j � r r f i l   ' % s ' .  K a n   i n t e   � p p n a   f j � r r f i l   ' % s ' .  K a n   i n t e   s t � n g a   f j � r r f i l   ' % s ' .  ' % s '   � r   i n t e   e n   f i l ! � � v e r f � r i n g e n   l y c k a d e s   s l u t f � r a ,   m e n   t e m p o r � r   � v e r f � r i n g s f i l   ' % s '   k u n d e   i n t e   b y t a   n a m n   t i l l   m � l f i l   ' % s ' .   O m   p r o b l e m e t   k v a r s t � r ,   p r o v a   m e d   a t t   s l �   a v   f i l � v e r f � r i n g e n s   � t e r u p p t a - f u n k t i o n  K a n   i n t e   s k a p a   l � n k   ' % s ' .  O g i l t i g t   k o m m a n d o   ' % s ' .  I n g e n 4 ' % s '   � r   i n g e n   t i l l � t e n   f i l r � t t i g h e t   i   o k t a l t   f o r m a t . 5 S e r v e r n   k r � v e r   e t t   e j   s t � t t   s l u t - p � - r a d   s e k v e n s   ( % s ) .  O k � n d   f i l t y p   ( % d )  O g i l t i g t   v e r k t y g .   % S � k v � g e n   f i n n s   i n t e   e l l e r   � r   o g i l t i g .  F i l e n   f i n n s   r e d a n . R F i l e n   l i g g e r   p �   e n   e n h e t   s o m   e n d a s t   s t � d e r   l � s n i n g ,   e l l e r   e n h e t e n   � r   s k r i v s k y d d a d .   D e t   f i n n s   i n g e t   m e d i a   i   e n h e t e n . * F e l   u p p s t o d   v i d   a v k o d n i n g   a v   U T F - 8   s t r � n g . < F e l   u p p s t o d   v i d   k � r n i n g   a v   e g e t   k o m m a n d o   ' % s '   p �   f i l e n   ' % s ' .  K a n   i n t e   l a d d a   l o c a l e   % d . + M o t t o g   e j   k o m p l e t t a   d a t a p a k e t   f � r e   f i l s l u t . 8 F e l   u p p s t o d   v i d   b e r � k n i n g   a v   s t o r l e k   f � r   k a t a l o g e n   ' % s ' . L M o t t o g   e t t   f � r   s t o r t   ( % d   B )   S F T P   p a k e t .   M a x i m a l t   s t � d d   p a k e t s t o r l e k   � r   % d   B . � K a n   i n t e   k � r a   S C P   f � r   a t t   s t a r t a   � v e r f � r i n g .   K o n t r o l l e r a   a t t   S C P   � r   i n s t a l l e r a t   p �   s e r v e r n   o c h   a t t   s � k v � g e n   � r   i n k l u d e r a d   i   P A T H .   D u   k a n   o c k s �   p r o v a   S F T P   i s t � l l e t   f � r   S C P .  P l a t s p r o f i l e n   ' % s '   f i n n s   r e d a n . , F e l   u p p s t o d   v i d   f l y t t   a v   f i l   ' % s '   t i l l   ' % s ' . x % s 
   
 F e l e t   o r s a k a s   n o r m a l t   a v   e t t   m e d d e l a n d e   f r � n   e t t   i n l o g g n i n g s s k r i p t   ( s o m   . p r o f i l e ) .   M e d d e l a n d e t   k a n   s t a r t a   m e d   " % s " . � U p p l a d d n i n g   a v   f i l e n   ' % s '   l y c k a d e s ,   m e n   e t t   f e l   u p p s t o d   n � r   f i l r � t t i g h e t e r n a   o c h / e l l e r   t i d s s t � m p e l n   s k u l l e   s � t t a s .   O m   p r o b l e m e t   k v a r s t � r ,   s l �   p �   a l t e r n a t i v e t   ' I g n o r e r a   r � t t i g h e t s f e l ' .  F e l a k t i g   m i n n e s � t k o m s t 2 D e t   f i n n s   i n g e n   l e d i g t   u t r y m m e   k v a r   i   f i l s y s t e m e t . t O p e r a t i o n e n   k a n   i n t e   s l u t f � r a s   p �   g r u n d   a v   a t t   d e t   s k u l l e   m e d f � r a   a t t   a n v � n d a r e n s   l a g r i n g s - q u o t a   s k u l l e   � v e r s k r i d a s . $ P r i n c i p a l   ( % s )   � r   o k � n t   f � r   s e r v e r n . 0 F e l   u p p s t o d   v i d   k o p i e r i n g   a v   f i l   ' % s '   t i l l   ' % s ' . ( O a v s l u t a t   m � n s t e r   ' % s '   v i d   b � r j a n   a v   % d . $ O k � n t   m � n s t e r   ' % s '   v i d   b � r j a n   a v   % d . V K a n   i n t e   k o m b i n e r a   f i l n a m n s m � n s t e r   ( b � r j a r   v i d   % d )   m e d   f i l l i s t m � n s t e r   ( b � r j a r   v i d   % d ) .  O k � n t   k o m m a n d o   ' % s ' . 0 T v e t y d i g t   k o m m a n d o   ' % s ' .   M � j l i g   m a t c h n i n g   � r :   % s $ P a r a m e t e r   s a k n a s   f � r   k o m m a n d o t   ' % s ' . ( F � r   m � n g a   p a r a m e t r a r   f � r   k o m m a n d o t   ' % s ' .  S e s s i o n e n   ' % s '   f i n n s   i n t e .        I n g e n   s e s s i o n .  O g i l t i g t   s e s s i o n s n u m m e r   ' % s ' .  O k � n t   a l t e r n a t i v   ' % s ' . % O k � n t   v � r d e   ' % s '   f � r   a l t e r n a t i v   ' % s ' . ( K a n   i n t e   b e s t � m m a   s t a t u s   p �   s o c k e t   ( % d ) . � F e l   u p p s t o d   v i d   b o r t t a g n i n g   a v   f i l   ' % s ' .   E f t e r   � t e r u p p t a g e n   f i l u p p l a d d n i n g   m � s t e   b e f i n t l i g   d e s t i n a t i o n s f i l   t a s   b o r t .   O m   d u   i n t e   h a   r � t t i g h e t e r   a t   t a   b o r t   d e s t i n a t i o n f i l ,   m � s t e   d u   a v a k t i v e r a   � t e r u p p t a g n i n g   a v   f i l � v e r f � r i n g . 5 F e l   u p p s t o d   v i d   a v k o d n i n g   a v   S F T P   p a k e t   ( % d ,   % d ,   % d ) . 1 O g i l t i g t   n a m n   ' % s ' .   N a m n   k a n   i n t e   i n n e h � l l a   ' % s ' . @ F i l e n   k u n d e   i n t e   � p p n a s   f � r   a t t   d e n   � r   l � s t   a v   e n   a n n a n   p r o c e s s .  K a t a l o g e n   � r   i n t e   t o m . + D e n   s p e c i f i c e r a d e   f i l e n   � r   i n t e   e n   k a t a l o g .  F i l n a m n e t   � r   i n t e   g i l t i g t . ( F � r   m � n g a   s y m b o l i s k a   l � n k a r   a n t r � f f a d e s .  F i l e n   k a n   i n t e   t a s   b o r t . p E n   a v   p a r a m e t r a r n a   v a r   u t a n f � r   i n t e r v a l l e t ,   e l l e r   p a r a m e t r a r n a   s o m   s p e c i f i c e r a d e s   k a n   i n t e   a n v � n d a s   t i l l s a m m a n s . V D e n   s p e c i f i c e r a d e   f i l e n   v a r   e n   k a t a l o g ,   i   e n   k o n t e x t   d � r   e n   k a t a l o g   i n t e   k a n   a n v � n d a s .  L � s   f � r   b y t e i n t e r v a l l   k r o c k a d e .  L � s   f � r   b y t e i n t e r v a l l   n e k a d e s . P E n   o p e r a t i o n   f � r s � k t e   g � r a s   p �   e n   f i l   s o m   h a r   e n   v � n t a n d e   b o r t t a g n i n g s o p e r a t i o n . F F i l e n   � r   k o r r u p t ;   e n   k o n t r o l l   a v   i n t e g r i t e t e n   i   f i l s y s t e m e t   b � r   k � r a s . L F i l e n   ' % s '   f i n n s   i n t e   e l l e r   d e n   i n n e h � l l e r   i n t e   p r i v a t   n y c k e l   i   k � n t   f o r m a t . � P r i v a t   n y c k e l f i l   ' % s '   i n n e h � l l e r   n y c k e l   i   % s   f o r m a t .   W i n S C P   s t � d e r   b a r a   P u T T Y   f o r m a t . 
   
 D u   k a n   a n v � n d a   P u T T Y g e n   v e r k t y g e t   f � r   a t t   k o n v e r t e r a   d i n   p r i v a t a   n y c k e l f i l . i P r i v a t   n y c k e l f i l   ' % s '   i n n e h � l l e r   n y c k e l   i   % s   f o r m a t .   D e n   f � l j e r   i n t e   d i n   f � r e d r a g n a   S S H   p r o t o k o l l v e r s i o n . z K a n   i n t e   s k r i v a   � v e r   f j � r r f i l   ' % s ' . 
   
 T r y c k   ' D e l e t e '   f � r   a t t   t a   b o r t   f i l   o c h   s k a p a   e n   n y   i s t � l l e t   f � r   a t t   s k r i v a   � v e r   d e n .  & T a   b o r t = F e l   u p p s t o d   v i d   k o n t r o l l   a v   l e d i g t   u t r y m m e   f � r   s � k v � g e n   ' % s ' . S K a n   i n t e   h i t t a   l e d i g   l o k a l   l i s t n i n g s p o r t n u m m e r   f � r   t u n n e l   i   i n t e r v a l l e t   % d   t i l l   % d . * K a n   i n t e   u t f � r a   n � t v e r k s h � n d e l s e   ( f e l   % d ) . / S e r v e r n   a v s l u t a d e   o v � n t a t   n � t v e r k s a n s l u t n i n g e n . 1 F e l   u p p s t o d   n � r   a n s l u t n i n g e n   s k u l l e   t u n n l a s . 
   
 % s 8 F e l   u p p s t o d   n � r   k o t r o l l s u m m a n   b e r � k n a d e s   f � r   f i l e n   ' % s ' .  I n t e r n t   f e l   % s   ( % s ) .  O p e r a t i o n e n   s t � d s   i n t e .    � t k o m s t   n e k a d .  F r � g a r   e f t e r   r e f e r e n s e r . . . $ O g i l t i g   s v a r   t i l l   P W D   k o m m a n d o   ' % s ' . + T h i s   v e r s i o n   d o e s   n o t   s u p p o r t   F T P   p r o t o c o l .  O k � n d   v � x e l   ' % s ' . ) F e l   u p p s t o d   v i d   � v e r f � r i n g   a v   f i l e n   ' % s ' .  K a n   i n t e   k � r a   ' % s ' .  F i l e n   ' % s '   h i t t a d e s   i n t e . . E t t   f e l   u p p s t o d   n � r   d o k u m e n t e t   s k u l l e   s t � n g a s . % ' % s '   � r   i n g e n   g i l t i g   h a s t i g h e t s g r � n s .              S j � l v s i g n e r a t   c e r t i f i k a t . , F o r m a t   f e l   i   c e r t i f i k a t e t s   g i l t i g - t i l l   f � l t . , F o r m a t   f e l   i   c e r t i f i k a t e t s   g i l t i g - f r � n   f � l t .  O g i l t i g   C A   c e r t i f i k a t .  E j   s t � t t   c e r t i f i k a t   � n d a m � l . 5 N y c k e l a n v � n d n i n g   i n k l u d e r a r   i n t e   c e r t i f i k a t s i g n e r i n g . , B e g r � n s n i n g a r   f � r   s � k v � g s l � n g d e n   � v e r s k r i d s . + S j � l v s i g n e r a t   c e r t i f i k a t   i   c e r t i f i k a t k e d j a . 6 D e t   g � r   i n t e   a t t   a v k o d a   u t f � r d a r e n s   o f f e n t l i g a   n y c k e l . 3 D e t   g � r   i n t e   a t t   d e k r y p t e r a   c e r t i f i k a t e t s   s i g n a t u r . ' D e t   g � r   i n t e   a t t   f �   u t f � r d a r c e r t i f i k a t . 2 D e t   g � r   i n t e   a t t   h � m t a   l o k a l t   u t f � r d a t   c e r t i f i k a t . 3 D e t   g � r   i n t e   a t t   v e r i f i e r a   d e t   f � r s t a   c e r t i f i k a t e t . % O k � n t   f e l   v i d   k o n t r o l l   a v   c e r t i f i k a t . 6 F e l e t   i n t r � f f a d e   p �   e t t   d j u p   a v   % d   i   c e r t i f i k a t k e d j a n .   C e r t i f i k a t e t   v e r k a r   v a r a   g i l t i g .    M a s k e n   � r   o g i l t i g   n � r a   ' % s ' . r S e r v e r n   k a n   i n t e   � p p n a   a n s l u t n i n g   i   a k t i v t   l � g e .   O m   p r o b l e m e t   k v a r s t � r ,   b � r   d u   � v e r v � g a   t t   b y t a   t i l l   p a s s i v t   l � g e . ( F e l   u p p s t o d   v i d   b o r t t a g n i n g   a v   f i l   ' % s ' .                    C O R E _ C O N F I R M A T I O N M V � r d e n   k o m m u n i c e r a r   i n t e   u n d e r   % d   s e k u n d e r . 
 
 V � n t a   y t t e r l i g a r e   % 0 : d   s e k u n d e r ?    & L � s e n o r d   f � r   n y c k e l n   ' % s ' :   # F i l e n   ' % s '   f i n n s   r e d a n .   S k r i v   � v e r ? ' K a t a l o g e n   ' % s '   f i n n s   r e d a n .   S k r i v   � v e r ? � D e t   f � r s t a   % s s k i f f r e t   s o m   s t � d s   a v   s e r v e r n   � r   % s ,   s o m   l i g g e r   u n d e r   k o n f i g u r e r a d   v a r n i n g s t r � s k e l n . 
 
 V i l l   d u   f o r t s � t t a   m e d   d e n   h � r   a n s l u t n i n g e n ?    k l i e n t - t i l l - s e r v e r  s e r v e r - t i l l - k l i e n t � M � l k a t a l o g e n   i n n e h � l l e r   d e n   d e l v i s   � v e r f � r d a   f i l e n   ' % s ' .   V i l l   d u   � t e r u p p t a   f i l � v e r f � r i n g e n ?   N o t e r a :   S v a r a s   ' N e j '   k o m m e r   a t t   t a   b o r t   d e n   d e l v i s   � v e r f � r d a   f i l e n   o c h   s t a r t a   � v e r f � r i n g e n   f r � n   b � r j a n . o M � l k a t a l o g e n   i n n e h � l l e r   d e n   d e l v i s   � v e r f � r d a   f i l e n   ' % s ' ,   s o m   � r   s t � r r e   � n   k � l l f i l e n .   F i l e n   k o m m e r   a t t   t a s   b o r t . y V i l l   d u   l � g g a   t i l l   f i l e n   ' % s '   t i l l   s l u t e t   p �   d e n   b e f i n t l i g a   f i l e n ?   V � l j   ' N e j '   f � r   a t t   � t e r u p p t a   f i l � v e r f � r i n g e n   i s t � l l e t . 4 % s 
   
 N y :             	 % s   b y t e s ,   % s 
 B e f i n t l i g :   	 % s   b y t e s ,   % s ' F i l e n   ' % s '   � r   s k r i v s k y d d a d .   S k r i v   � v e r ? ' L o k a l   f i l   ' % s '   f i n n s   r e d a n .   S k r i v   � v e r ? & F j � r r f i l   ' % s '   f i n n s   r e d a n .   S k r i v   � v e r ?           C V � r d e n   k o m m u n i c e r a r   i n t e   p �   � v e r   % d   s e k u n d e r .   V � n t a r   f o r t f a r a n d e . . . � D e n   f � r s t a   a l g o r i t m e n   f � r   n y c k e l u t b y t e   s o m   s t � d s   a v   s e r v e r n   � r   % s ,   s o m   l i g g e r   u n d e r   k o n f i g u r e r a d   v a r n i n g s t r � s k e l . 
 
 V i l l   d u   f o r t s � t t a   m e d   d e n   h � r   a n s l u t n i n g e n ?  & � t e r a n s l u t 
 N y t t   n a & m n      T u n n e l   f � r   % s  L � s e n o r d  L � s e n o r d   f � r   n y c k e l  S e r v e r p r o m p t  A n v � n d a r n a m n  A & n v � n d a r n a m n :  S e r v e r p r o m p t :   % s  N y t t   l � s e n o r d  S & v a r :    A n v � n d e r   T I S   a u t e n t i s e r i n g . % s $ A n v � n d e r   K r y p t o k o r t   a u t e n t i s e r i n g . % s 
 & L � s e n o r d : / A n v � n d e r   t a g e n t b o r d s i n t e r a k t i v   a u t e n t i s e r i n g . % s  N & u v a r a n d e   l � s e n o r d :  & N y t t   l � s e n o r d  & B e k r � f t a   n y t t   l � s e n o r d :  A u t e n t i s e r i n g   f � r   t u n n e l s e s s i o n  � v e r f � r   m e d   e t t   a n n a t   n a m n  & N y t t   n a m n : TS e r v e r n s   c e r t i f i k a t   � r   i n t e   k � n t .   D u   h a r   i n g e n   g a r a n t i   a t t   s e r v e r n   � r   d e n   d a t o r n   d u   t r o r   d e t   � r .   S e r v e r n s   c e r t i f i k a t i n f o r m a t i o n   f � l j e r : 
 
 % s 
 
 O m   d u   l i t a r   p �   d e t   h � r   c e r t i f i k a t e t ,   t r y c k   p �   J a .   O m   d u   v i l l   a n s l u t a   u t a n   a t t   s p a r a   c e r t i f i k a t e t ,   t r y c k   p �   N e j .   F � r   a t t   � v e r g e   a n s l u t n i n g e n ,   t r y c k   p �   A v b r y t . 
 
 F o r t s � t t   a n s l u t a   o c h   l a g r a   c e r t i f i k a t e t ? - -   O r g a n i s a t i o n :   % s 
 | -   P l a t s :   % s 
 | -   A n n a t :   % s 
  % s ,   % s S U t g i v a r e : 
 % s 
 � m n e : 
 % s 
 G i l t i g :   % s   -   % s 
 
 F i n g e r a v t r y c k   ( S H A 1 ) :   % s 
 
 S a m m a n f a t t n i n g :   % s      C O R E _ I N F O R M A T I O N  J a  N e j ` V � r d :   % s 
 A n v � n d a r n a m n :   % s 
 P r i v a t   n y c k e l f i l :   % s 
 S S H   p r o t o k o l l v e r s i o n :   % s 
 � v e r f � r i n g s p r o t o k o l l :   % s  V e r s i o n   % d . % d . % d   ( B y g g d   % d ) > O p e r a t i o n e n   s l u t f � r d e s   f r a m g � n g s r i k t .   A n s l u t n i n g e n   a v s l u t a d e s .  S F T P - % d : S F T P   p r o t o k o l l e t s   v e r s i o n   t i l l � t e r   i n t e   n a m n b y t e   p �   f i l e r . ' S e r v e r n   s t � d e r   i n g a   u t � k n i n g a r   a v   S F T P . ( S e r v e r n   s t � d e r   f � l j a n d e   S F T P   u t � k n i n g a r :     
 L � & g g   t i l l  E n d a s t   n & y a r e  V i s a r   h j � l p . S t � n g e r   a l l a   s e s s i o n e r   o c h   a v s l u t a r   p r o g r a m m e t  A n s l u t e r   t i l l   s e r v e r  S t � n g e r   s e s s i o n e n 4 L i s t a r   a n s l u t n a   s e s s i o n e r   e l l e r   v � l j e r   a k t i v   s e s s i o n  V i s a r   a k t u e l l   f j � r r k a t a l o g  B y t e r   a k t u e l l   f j � r r k a t a l o g  V i s a r   i n n e h � l l e t   i   f j � r r k a t a l o g  V i s a r   a k t u e l l   l o k a l   k a t a l o g  B y t e r   a k t u e l l   l o k a l   k a t a l o g ! L i s t a r   i n n e h � l l e t   i   l o k a l   k a t a l o g  T a r   b o r t   f j � r r f i l  T a r   b o r t   f j � r r k a t a l o g $ F l y t t a r   e l l e r   b y t e r   n a m n   p �   f j � r r f i l   � n d r a r   r � t t i g h e t e r n a   p �   f j � r r f i l  S k a p a r   e n   s y m b o l i s k   f j � r r l � n k  S k a p a r   f j � r r k a t a l o g 3 L a d d a r   n e r   f i l   f r � n   f j � r r k a t a l o g   t i l l   l o k a l   k a t a l o g 3 L a d d a r   u p p   f i l   f r � n   l o k a l   k a t a l o g   t i l l   f j � r r k a t a l o g - S � t t e r   e l l e r   v i s a r   v � r d e n   p �   s c r i p t a l t e r n a t i v , S y n k r o n i s e r a r   f j � r r k a t a l o g   m e d   l o k a l   k a t a l o g D K o n t i n u e r l i g t   � t e r s p e g l a   � n d r i n g a r   i   l o k a l   k a t a l o g   t i l l   f j � r r k a t a l o g  V � r d :      A k t i v   s e s s i o n :   [ % d ]   % s  S e s s i o n   ' % s '   a v s l u t a d .  L o k a l   ' % s '   % s   F j � r r   ' % s '  ' % s '   b o r t t a g e n 7 � v e r v a k a r   f � r � n d r i n g a r ,   t r y c k   C T R L - C   f � r   a t t   a v b r y t a . . .  & H o p p a   � v e r   a l l a  K � r   g o d t y c k l i g t   f j � r r k o m m a n d o  & T e x t  & B i n � r t  & U t e s l u t   t i l l f � l l i g a / � v e r f � r i n g s t y p :   % s | B i n � r t | T e x t | A u t o m a t i s k t   ( % s ) O F i l n a m n s f � r � n d r i n g :   % s | I n g e n   � n d r i n g | V e r s a l e r | G e m e n e r | F � r s t a   v e r s a l | G e m e n e r   8 . 3  S � t t   r � t t i g h e t e r :   % s  L � g g   t i l l   X   t i l l   k a t a l o g  B e v a r a   t i d s s t � m p e l  U t e s l u t   m a s k :   % s  I n k l u d e r a   m a s k :   % s  R e n s a   ' A r k i v '   a t t r i b u t  B y t   i n t e   u t   o g i l t i g a   t e c k e n    B e v a r a   i n t e   t i d s s t � m p e l  B e r � k n a   i n t e   � v e r f � r i n g s s t o r l e k   S t a n d a r d � v e r f � r i n g s i n s t � l l n i n g a r  V � r d n a m n :   % s  A n v � n d a r n a m n :   % s  F j � r r k a t a l o g :   % s    L o k a l   k a t a l o g :   % s $ S k a n n a r   ' % s '   e f t e r   u n d e r k a t a l o g e r . . . % � v e r v a k a r   � n d r i n g a r   i   % d   k a t a l o g e r . . .  � n d r i n g   i   ' % s '   u p p t � c k t .  F i l   ' % s '   u p p l a d d a d .  F i l   ' % s '   b o r t t a g e n . U % s   k o n f i g u r e r a d   � v e r f � r i n g s i n s t � l l n i n g   k a n   i n t e   a n v � n d a s   i   a k t u e l l   k o n t e x t | N � g o n | A l l a    I g n o r e r a   r � t t i g h e t s f e l  A n v � n d e r   a n v � n d a r n a m n   " % s " . . A n v � n d e r   t a n g e n t b o r d s i n t e r a k t i v   a u t e n t i s e r i n g . % A u t e n t i s e r i n g   m e d   p u b l i k   n y c k e l   " % s " .  F e l a k t i g   l � s e n o r d .  � t k o m s t   n e k a d . 0 A u t e n t i s e r i n g   m e d   p u b l i k   n y c k e l   " % s "   f r � n   a g e n t . ( F � r s � k e r   m e d   p u b l i k   n y c k e l a u t e n t i s e r i n g .   ' A u t e n t i s e r i n g   m e d   f � r i n s t � l l t   l � s e n o r d .  � p p n a r   t u n n e l . . .  A n s l u t n i n g   a v s l u t a d .    S � k e r   e f t e r   v � r d . . .  A n s l u t e r   t i l l   v � r d . . .  A u t e n t i s e r a r . . .  A u t e n t i s e r a d .  S t a r t a r   s e s s i o n e n . . .  L � s e r   f j � r r k a t a l o g . . .  S e s s i o n e n   s t a r t a d .  A n s l u t e r   g e n o m   t u n n e l . . .  S e r v e r   n e k a r   v � r   n y c k e l .  A d m i n i s t r a t i v t   f � r b j u d e n   ( % s ) .  A n s l u t n i n g   m i s s l y c k a d e s   ( % s ) .  N � t v e r k s f e l :   A n s l u t n i n g   n e k a s .   + N � t v e r k s f e l :   A n s l u t n i n g   � t e r s t � l l d   a v   p e e r .   N � t v e r k s f e l :   A n s l u t n i n g s t i m e o u t . 2 V � r d :   % s 
 A n v � n d a r n a m n :   % s 
 � v e r f � r i n g s p r o t o k o l l :   % s 
 & � t e r u p p t a / S e r v e r n   s t � d e r   i n t e   n � g r a   e x t r a   F T P   e g e n s k a p e r . . S e r v e r n   s t � d e r   d e   h � r   e x t r a   F T P   e g e n s k a p e r n a :   $ � v e r f � r i n g s h a s t i g h e t s g r � n s :   % u   K i B / s  & K o p i e r a   n y c k e l 
 & U p p d a t e r a 
 & L � g g   t i l l  B e v a r a   e n d a s t   l � s n i n g 	 J � m f � r . . .  S y n k r o n i s e r a r . . .  I n g e t   a t t   s y n k r o n i s e r a . 
 O b e g r � n s a d  S S L / T L S   I m p l i c i t   k r y p t e r i n g    S S L   E x p l i c i t   k r y p t e r i n g  T L S   E x p l i c i t   k r y p t e r i n g                                              C O R E _ V A R I A B L E ( S S H   o c h   S C P   k o d e n   � r   b a s e r a d   p �   P u T T Y   % s  0 . 6 0 " C o p y r i g h t   �   1 9 9 7 - 2 0 0 9   S i m o n   T a t h a m 2 h t t p : / / w w w . c h i a r k . g r e e n e n d . o r g . u k / ~ s g t a t h a m / p u t t y / $ F T P   k o d e n   � r   b a s e r a d   p �   F i l e Z i l l a   % s  2 . 2 . 3 2  C o p y r i g h t   �   2 0 0 1 - 2 0 0 7   T i m   K o s s e ! h t t p : / / f i l e z i l l a . s o u r c e f o r g e . n e t / m D e n n a   p r o d u k t   i n n e h � l l e r   p r o g r a m v a r a   s o m   u t v e c k l a t s   a v   O p e n S S L   P r o j e c t   f � r   a n v � n d n i n g   i   O p e n S S L : s   v e r k t y g   % s . ) C o p y r i g h t   �   1 9 9 8 - 2 0 0 9   T h e   O p e n S S L   P r o j e c t  0 . 9 . 8 k  h t t p : / / w w w . o p e n s s l . o r g /                                           �D u   f � r s � k e r   f l y t t a   f j � r r f i l e r   t i l l   e n   d e s t i n a t i o n   s o m   W i n S C P   i n t e   k a n   f l y t t a   t i l l   d i r e k t .   F i l e r n a   k o m m e r   a t t   l a d d a s   n e r   t i l l   e n   t e m p o r � r   k a t a l o g   i s t � l l e t .   A n s v a r e t   f � r   � v e r f � r i n g e n   t i l l   d e n   s l u t g i l t i g a   d e s t i n a t i o n e n   s k a   s k � t a s   a v   m � l a p p l i k a t i o n e n   ( t .   e x .   U t f o r s k a r e n ) ,   v i l k e t   W i n S C P   i n t e   k a n   k o n t r o l l e r a .   K � l l f i l e r   k o m m e r   a t t   r a d e r a s   e f t e r   a t t   n e r l a d d n i n g e n   t i l l   d e n   t e m p o r � r a   k a t a l o g e n   h a r   a v s l u t a t s .   O m   m � l a p p l i k a t i o n e n   m i s s l y c k a s   m e d   a t t   h a n t e r a   d e   t e m p o r � r a   f i l e r n a ,   k a n   d e   f � r l o r a s .   � v e r v � g   g � r n a   a t t   k o p i e r a   f i l e r n a   i s t � l l e t   f � r   a t t   f l y t t a   d e m . 
 T i p s :   F � r   a t t   k o p i e r a   f i l e r   h � l l   n e r   C T R L   t a n g e n t e n   m e d a n   f l y t t . 
 
 V i l l   d u   f o r t f a r a n d e   f l y t t a   f i l e r n a ? YW i n S C P ,   % s 
 % s 
 
 A n v � n d n i n g : 
 G : % A P P %   s e s s i o n 
 G : % A P P %   [ ( s f t p | s c p | f t p ) : / / ] [ u s e r [ : p a s s w o r d ] @ ] h o s t [ : p o r t ] [ / p a t h / [ f i l e ] ] 
 G : % A P P %   [ s e s s i o n ]   / s y n c h r o n i z e   [ l o c a l _ d i r ]   [ r e m o t e _ d i r ]   [ / d e f a u l t s ] 
 G : % A P P %   [ s e s s i o n ]   / k e e p u p t o d a t e   [ l o c a l _ d i r ]   [ r e m o t e _ d i r ]   [ / d e f a u l t s ] 
 G : % A P P %   [ s e s s i o n ]   / p r i v a t e k e y = < k e y >   / h o s t k e y = < f i n g e r p r i n t > 
 G : % A P P %   [ s e s s i o n ]   / c e r t i f i c a t e = < f i n g e r p r i n t >   / i m p l i c i t | e x p l i c i t s s l | e x p l i c i t t l s 
 G : % A P P %   [ s e s s i o n ]   / p a s s i v e   / t i m e o u t = < s e c > 
 G : % A P P %   [ / c o n s o l e ]   [ / s c r i p t = f i l e ]   [ / c o m m a n d   c o m m a n d 1 . . . ]   [ / p a r a m e t e r   p a r a m 1 . . . ] 
 C : % A P P %   [ / s c r i p t = f i l e ]   [ / c o m m a n d   c o m m a n d 1 . . . ]   [ / p a r a m e t e r   p a r a m 1 . . . ] 
 B : % A P P %   / i n i = < i n i f i l e >   / l o g = < l o g f i l e > 
 G : % A P P %   / u p d a t e 
 B : % A P P %   / h e l p 
 
 G :   s e s s i o n               N a m n   p �   l a g r a d   s e s s i o n   e l l e r   d i r e k t   s e s s i o n s s p e c i f i k a t i o n . 
 G :   / s y n c h r o n i z e     S y n k r o n i s e r a r   i n n e h � l l e t   i   t v �   k a t a l o g e r . 
 G :   / k e e p u p t o d a t e   S t a r t a r   f u n k t i o n e n :   H � l l   f j � r r k a t a l o g e n   a k t u e l l . 
 G :   / d e f a u l t s           S t a r t a r   o p e r a t i o n e n   u t a n   a t t   v i s a   d i a l o g r u t a n   A l t e r n a t i v . 
 G :   / c o n s o l e             K o n s o l l   ( t e x t )   - l � g e .   S t a n d a r d l � g e t ,   n � r   d e n   a n r o p a s 
 G :                               g e n o m   % A P P % . c o m . 
 B :   / s c r i p t =             K � r   b a t c h - s k r i p t f i l .   O m   i n t e   s k r i p t e t   s l u t a r   m e d 
 B :                               ' e x i t '   k o m m a n d o ,   n o r m a l t   i n t e r a k t i v t   l � g e   f � l j e r . 
 B :   / c o m m a n d             K � r   l i s t a   � v e r   s k r i p t k o m m a n d o n . 
 B :   / p a r a m e t e r         S k i c k a r   l i s t a   m e d   p a r a m e t r a r   t i l l   s k r i p t . 
 B :   / i n i =                   S � k v � g   t i l l   k o n f i g u r a t i o n s   I N I - f i l . 
 B :   / l o g =                   S t a r t a r   l o g g n i n g   t i l l   f i l . 
 G :   / p r i v a t e k e y =     P r i v a t   n y c k e l f i l . 
 G :   / t i m e o u t =           S e r v e r s v a r   t i m e o u t . 
 G :   / h o s t k e y =           F i n g e r a v t r y c k   f � r   s e r v e r n s   v � r d n y c k e l . 
 G :   / p a s s i v e             P a s s i v t   l � g e   ( e n d a s t   F T P   p r o t o k o l l ) . 
 G :   / c e r t i f i c a t e =   F i n g e r a v t r y c k   f � r   S S L / T L S   c e r t i f i k a t . 
 G :   / i m p l i c i t           I m p l i c i t   T L S / S S L   ( e n d a s t   F T P S   p r o t o k o l l ) . 
 G :   / e x p l i c i t s s l     E x p l i c i t   S S L   ( e n d a s t   F T P S   p r o t o k o l l ) . 
 G :   / e x p l i c i t t l s     E x p l i c i t   T L S   ( e n d a s t   F T P S   p r o t o k o l l ) . 
 G :   / u p d a t e               F r � g a r   a p p l i k a t i o n e n s   h e m s i d a   o m   u p p d a t e r i n g a r . 
 B :   / h e l p                   S k r i v e r   d e n n a   a n v � n d n i n g . 
                                   	 W I N _ E R R O R   Q % s 
   
 V a r n i n g :   A t t   a v b r y t a   d e n   h � r   o p e r a t i o n e n   k o m m e r   a t t   s t � n g a   n e r   a n s l u t n i n g e n !          K a n   i n t e   s k a p a   g e n v � g . ) K a n   i n t e   s k r i v a   � v e r   s p e c i a l s e s s i o n   ' % s ' .  K a n   i n t e   u t f o r s k a   k a t a l o g   ' % s ' . , I n g e n   f i l l i s t a   f � r   u p p l a d d n i n g   h a r   a n g i v i t s .  K a n   i n t e   s k a p a   m a p p e n   ' % s ' .   ' K a n   i n t e   t a   b o r t   t e m p o r � r   k a t a l o g   ' % s ' . % K a n   i n t e   � p p n a   e l l e r   k � r a   f i l e n   ' % s ' .  K a n   i n t e   s t a r t a   e d i t o r   ' % s ' .   w K a n   i n t e   � p p n a   m o t s v a r a d e   k a t a l o g   i   m o t s a t t   p a n e l .   S y n k r o n i s e r i n g   a v   k a t a l o g b l � d d r i n g   m i s s l y c k a d e s .   D e n   h a r   s t � n g t s   a v .  K a n   i n t e   a v g � r a   g e n v � g   ' % s ' .   % ' % s '   � r   i n t e   g i l t i g t   p l a t s p r o f i l n a m n . 1 ' % s '   � r   i n t e   g i l t i g t   n a m n   f � r   e n   p l a t s p r o f i l m a p p . , P l a t s p r o f i l m a p p   m e d   n a m n e t   ' % s '   f i n n s   r e d a n . 5 B e s k r i v n i n g   p �   e g e t   k o m m a n d o   k a n   i n t e   i n n e h � l l a   ' % s ' . 1 E g e t   k o m m a n d o   m e d   b e s k r i v n i n g e n   ' % s '   f i n n s   r e d a n . D K a n   i n t e   f r � g a   a p p l i k a t i o n e n s   h e m s i d a   e f t e r   u p p d a t e r i n g s i n f o r m a t i o n . , F e l   u p p s t o d   v i d   s � k n i n g   e f t e r   u p p d a t e r i n g a r .         P K a n   i n t e   r e g i s t r e r a   a p p l i k a t i o n e n   f � r   a t t   h a n t e r a   a d r e s s e r n a   s c p : / /   o c h   s f t p : / / . 2 M u t e x   s l � p p t e s   i n t e   e n l i g t   d e t   k r � v d a   i n t e r v a l l e t . E S k a l   d r a - t i l l � g g e t   m u t e x   s l � p p t e s   i n t e   e n l i g t   d e t   k r � v d a   i n t e r v a l l e t . �W i n S C P   k u n d e   i n t e   h i t t a   m a p p e n ,   d � r   d e   d r a g n a   f i l e r n a   s l � p p t e s .   A n t i n g e n   h a r   f i l e r n a   i n t e   s l � p p t s   t i l l   e n   v a n l i g   m a p p   ( t .   e x .   i   U t f o r s k a r e n )   e l l e r   s �   � r   W i n S C P   s k a l   d r a - t i l l � g g e t   i n t e   i n s t a l l e r a d   e l l e r   h a r   d u   i n t e   s t a r t a t   o m   d a t o r n   e f t e r   i n s t a l l a t i o n .   I n s t a l l e r a   t i l l � g g e t   e l l e r   v � l j   e t t   k o m p a t i b e l t   d r a   & &   s l � p p - l � g e   ( i   i n s t � l l n i n g s f � n s t r e t ) ,   s o m   a n v � n d e r   s i g   a v   e n   t e m p o r � r   m a p p   v i d   n e r l a d d n i n g .   D e t t a   m � j l i g g � r   a t t   d r a   f i l e r   t i l l   v a l f r i   d e s t i n a t i o n . K F i l e n   ' % s '   i n n e h � l l e r   i n t e   n � g o n   � v e r s � t t n i n g   f � r   d e n   h � r   p r o d u k t v e r s i o n e n . 5 F i l e n   ' % s '   i n n e h � l l e r   � v e r s � t t n i n g   f � r   % s   v e r s i o n   % s . 6S k a l e t s   d r a   & &   s l � p p - t i l l � g g   � r   p � s l a g e t ,   m e n   t i l l � g g e t   l a d d a d e s   i n t e .   A n t i n g e n   � r   t i l l � g g e t   i n t e   i n s t a l l e r a t   e l l e r   s �   h a r   d a t o r n   i n t e   s t a r t a t s   o m   e f t e r   i n s t a l l a t i o n e n .   I n s t a l l e r a   t i l l � g g e t   e l l e r   v � x l a   t i l l   e t t   k o m p a t i b e l t   d r a   & &   s l � p p - l � g e   ( v i a   I n s t � l l n i n g a r ) ,   s o m   a n v � n d e r   e n   t e m p o r � r   m a p p   f � r   n e r l a d d n i n g a r . 8 G S S A P I / S S P I   m e d   K e r b e r o s   s t � d s   i n t e   p �   d e t   h � r   s y s t e m e t . ' F e l   u p p s t o d   v i d   b e v a k n i n g   a v   � n d r i n g a r . 8 F e l   u p p s t o d   v i d   b e v a k n i n g   a v   � n d r i n g a r   i   k a t a l o g e n   ' % s ' .   6 F e l   u p p s t o d   v i d   b e v a k n i n g e n   a v   � n d r i n g a r   i   f i l e n   ' % s ' . L K a n   i n t e   l a d d a   u p p   r e d i g e r a d   f i l   ' % s ' ,   s e s s i o n e n   ' % s '   h a r   r e d a n   s t � n g t s   n e r . I D e t   f i n n s   r e d a n   f � r   m � n g a   f i l e r   � p p n a d e .   V a r   g o d   s t � n g   n � g r a   f i l e r   f � r s t .   R % s   V a r   v � n l i g   t a   b o r t   f i l e n .   A n n a r s   k o m m e r   i n t e   a p p l i k a t i o n e n   a t t   f u n g e r a   k o r r e k t . o K a n   i n t e   s k a p a   t e m p o r � r   k a t a l o g   ' % s ' .   D u   k a n   � n d r a   r o t k a t a l o g e n   f � r   l a g r i n g   a v   t e m p o r � r a   f i l e r   i   I n s t � l l n i n g a r . �W i n S C P   k u n d e   i n t e   a v g � r a   v i l k e t   p r o g r a m   s o m   s k a   s t a r t a s   f � r   a t t   � p p n a   f i l e n .   W i n S C P   k a n   i n t e   b e v a k a   � n d r i n g a r   i   f i l e n ,   s �   d e n   v i l l   i n t e   l a d d a s   u p p . 
   
 E n   m � j l i g   o r s a k   t i l l   p r o b l e m e t   � r   a t t   f i l e n   r e d a n   h a r   � p p n a t s   a v   e t t   a n n a t   p r o g r a m   s o m   k � r s . 
   
 O m   d u   v i l l   a n v � n d a   p r o g r a m m e t   f � r   a t t   � p p n a   f i l e r   f r � n   W i n S C P ,   � v e r v � g   a t t   k o n f i g u r e r a   d e n   s o m   e n   e x t e r n   e d i t o r . 
   
 N o t e r a   a t t   f i l e n   l i g g e r   k v a r   i   d e n   t e m p o r � r a   m a p p e n . � N � g r a   a v   d e   t e m p o r � r a   m a p p a r n a   k u n d e   i n t e   t a s   b o r t .   O m   f i l e r   f i n n s   l a g r a d e   d � r   s o m   f o r t f a r a n d e   � r   � p p n a ,   s t � n g   d e s s a   o c h   p r o v a   i g e n . � F � r   a t t   a n v � n d a   v a l t   e g e t   k o m m a n d o ,   f � r   b a r a   e n   f i l   v a r a   m a r k e r a d   i   d e n   e n a   p a n e l e n ,   f � r   a t t   k � r a   k o m m a n d o t   p �   d e   v a l d a   f i l e r n a   i   m o t s a t t   p a n e l .   A l t e r n a t i v t   k a n   s a m m a   a n t a l   f i l e r   m a r k e r a s   i   b � d a   p a n e l e r n a   f � r   a t t   k � r a   k o m m a n d o t   p �   m a t c h a n d e   p a r   a v   f i l e r . W F � r   a t t   a n v � n d a   v a l t   e g e t   k o m m a n d o t   f � r   b a r a   e n   f i l   v a r a   m a r k e r a d   i   d e n   l o k a l a   p a n e l e n .   � N � g r a   a v   d e   v a l d a   f j � r r f i l e r n a   l a d d a d e s   i n t e   n e r .   D e t   v a l d a   e g n a   k o m m a n d o t   m � s t e   k � r a s   p �   m a t c h a n d e   p a r   a v   f i l e r ,   v i l k e t   d � r f � r   i n t e   � r   m � j l i g t . $ K a n   i n t e   i n i t i a l i s e r a   e x t e r n   k o n s o l . C M e d d e l a n d e t   f � r   l � n g t   ( % d   b y t e s )   f � r   a t t   s k i c k a   t i l l   e x t e r n   k o n s o l . N K a n   i n t e   � p p n a   m a p p n i n g s o b j e k t   f � r   a t t   s t a r t a   k o m m u n i k a t i o n   m e d   e x t e r n   k o n s o l . ; T i m e o u t   v � n t a r   p �   e x t e r n   k o n s o l   f � r   a t t   s l u t f � r a   k o m m a n d o t . 4 I n k o m p a t i b e l t   p r o t o k o l l v e r s i o n   f � r   e x t e r n   k o n s o l   % d . E F e l   u p p s t o d   n � r   s � k v � g   ' % s '   l a d d e s   t i l l   m i l j � v a r i a b e l   p a t h ( % % P A T H % % ) . H F e l   u p p s t o d   n � r   s � k v � g   ' % s '   t o g s   b o r t   f r � n   m i l j � v a r i a b e l   p a t h ( % % P A T H % % ) .   [ F i l e n   ' % s '   � r   r e d a n   � p p n a d   i   e n   e x t e r n   e d i t o r   ( a p p l i k a t i o n )   e l l e r   h � l l e r   p �   a t t   l a d d a s   u p p . 8 D u   h a r   i n t e   a n g i v i t   n � g o n   a u t o m a t i s k t   v a l   a v   m a s k r e g l e r . D F � r i n s t � l l d   � v e r f � r i n g s i n s t � l l n i n g   m e d   b e s k r i v n i n g   ' % s '   f i n n s   r e d a n . K E g e t   k o m m a n d o   ' % s '   k a n   i n t e   k � r a s   j u s t   n u .   V � l j   f � r s t   f i l e r   t i l l   k o m m a n d o t . A K a n   i n t e   l a d d a   o m   f i l e n   ' % s ' ,   s e s s i o n e n   ' % s '   h a r   r e d a n   a v s l u t a t s .   S A u t o m a t i s k a   � t g � r d e r   � r   a v s t � n g d a   n � r   U R L   a d r e s s e n   t i l l h a n d a h � l l s   p �   k o m m a n d o r a d e n .     L � s e n o r d e t   k a n   i n t e   d e k r y p t e r a s . 3 D u   h a r   i n t e   a n g e t t   k o r r e k t   n u v a r a n d e   h u v u d l � s e n o r d . 0 N y a   o c h   u p p r e p a d e   h u v u d l � s e n o r d e t   � r   i n t e   s a m m a .                                      W I N _ C O N F I R M A T I O N . S e s s i o n   m e d   n a m n   ' % s '   f i n n s   r e d a n .   S k r i v   � v e r ? ! K a t a l o g e n   ' % s '   f i n n s   i n t e .   S k a p a ?  A v b r y t   a k t u e l l   o p e r a t i o n ? � A v b r y t   f i l � v e r f � r i n g ? 
   
 O p e r a t i o n e n   k a n   i n t e   a v b r y t a s   m i t t   u n d e r   f i l � v e r f � r i n g . 
 V � l j   ' J a '   f � r   a t t   a v b r y t a   f i l � v e r f � r i n g e n   o c h   s t � n g a   a n s l u t n i n g e n . 
 V � l j   ' N e j '   f � r   a t t   f u l l f � l j a   f i l � v e r f � r i n g e n . 
 V � l j   ' A v b r y t '   f � r   a t t   f o r t s � t t a   o p e r a t i o n e n . . � r   d u   s � k e r   p �   a t t   d u   v i l l   t a   b o r t   f i l e n   ' % s ' ? 7 � r   d u   s � k e r   p �   a t t   d u   v i l l   t a   b o r t   d e   % d   v a l d a   f i l e r n a ? / A v s l u t a   s e s s i o n e n   ' % s '   o c h   s t � n g   a p p l i k a t i o n e n ?  F r � g a   m i & g   a l d r i g   i g e n <F � r   l i t e   l e d i g t   u t r y m m e   p �   t e m p o r � r   e n h e t ! 
 
 N � r   f i l e r   d r a s   f r � n   e n   f j � r r k a t a l o g ,   l a d d a s   f i l e r n a   f � r s t   n e r   t i l l   e n   t e m p o r � r   k a t a l o g   ' % s ' .   D e t   � r   % s   l e d i g t   p �   e n h e t e n .   T o t a l   s t o r l e k   f � r   d e   v a l d a   f i l e r n a   � r   % s . 
 
 N o t e r a :   T e m p o r � r   k a t a l o g e n   k a n   � n d r a s   i   I n s t � l l n i n g s f � n s t r e t . 
 
 V i l l   d u   f o r t s � t t a   m e d   a t t   l a d d a   n e r   f i l e r n a ?   ( L � g g   t i l l   k a t a l o g e n   ' % s '   t i l l   b o k m � r k e n ?     - S k a p a   g e n v � g   p �   s k r i v b o r d e t   f � r   s e s s i o n   ' % s ' ? 2 A n v � n d   a k t u e l l a   s e s s i o n s i n t � l l n i n g a r   s o m   s t a n d a r d ?  & H o p p a   � v e r # F i l e n   h a r   � n d r a t s .   S p a r a   � n d r i n g a r ? 9 S k a p a   u t f o r s k a r e n s   ' S k i c k a   t i l l ' - g e n v � g   f � r   s e s s i o n   ' % s ' ?  S k a p a   v a l d   i k o n / g e n v � g ? / A v s l u t a   a l l a   s e s s i o n e r   o c h   s t � n g   a p p l i k a t i o n e n ?  T a   b o r t   v a l d   p l a t s p r o f i l m a p p ?  & F � r e g � e n d e  & N � s t a   V V i l l   d u   a t t   a p p l i k a t i o n e n   r e g i s t r e r a s   f � r   a t t   h a n t e r a   a d r e s s e r   m e d   s c p : / /   o c h   s f t p : / / ? L V i l l   d u   r e n s a   u p p   d a t a   f r � n   d e n   h � r   d a t o r n   s o m   h a r   s k a p a t s   a v   a p p l i k a t i o n e n ? ! % s 
 
 V i l l   d u   s t � n g a   a p p l i k a t i o n e n ? G % % s 
 
 V i l l   d u   a v s l u t a   % d   � t e r s t � e n d e   s e s s i o n e r   o c h   s t � n g a   a p p l i k a t i o n e n ? � D e t   f i n n s   f o r t f a r a n d e   b a k g r u n d s � v e r f � r i n g a r   i   k � n .   V i l l   d u   k o p p l a   i f r � n   � n d � ? 
   
 V a r n i n g :   A t t   v � l j a   ' O K '   k o m m e r   a t t   a v s l u t a   a l l a   p � g � e n d e   � v e r f � r i n g a r .  A k t u e l l   s e s s i o n   % s   s t � d e r   i n t e   d e t   a k t u e l l a   k o m m a n d o t .   E n   s e p a r a t   s k a l s e s s i o n   k o m m e r   a t t   � p p n a s   f � r   a t t   u t f � r a   k o m m a n d o t .   S k a   e n   s e p a r a t   s k a l s e s s i o n   � p p n a s ? 
   
 N o t e r a :   S e r v e r n   m � s t e   t i l l h a n d a h � l l a   e t t   U n i x - l i k n a n d e   s k a l   o c h   s k a l e t   m � s t e   a n v � n d a   s a m m a   s � k v � g s - s y n t a x   s o m   a k t u e l l   s e s s i o n   % s . � D e t   f i n n s   n � g r a   � p p n a   f i l e r .   V a r   v � n l i g   s t � n g   d e m   i n n a n   a p p l i k a t i o n e n   a v s l u t a s . 
   
 N o t e r a :   O m   d e t t a   i n t e   u t f � r s ,   k a n   r e d i g e r a d e   f i l e r   l i g g a   k v a r   i   d e n   t e m p o r � r a   k a t a l o g e n . W i n S C P   h i t t a d e   % d   t e m p o r � r a   m a p p a r ,   s o m   a n t a g l i g e n   h a r   s k a p a t s   t i d i g a r e .   D e s s a   m a p p a r   k a n   i n n e h � l l a   f i l e r   s o m   t i d i g a r e   h a r   r e d i g e r a t s   e l l e r   l a d d a t s   n e r .   V i l l   d u   t a   b o r t   d e s s a   m a p p a r ?   D u   k a n   o c k s �   � p p n a   m a p p a r n a   f � r   a t t   s e   i n n e h � l l e t   o c h   t a   b o r t   d e m   m a n u e l l t .  & � p p n a # V i s a   i n t e   d e t   h � r   m e d d e l a n d e t   i & g e n   ` V i l l   d u   s k a p a   s k r i v b o r d i k o n   f � r   a l l a   a n v � n d a r e ? 
   
 D u   m � s t e   h a   a d m i n i s t r a t � r s r � t t i g h e t e r   f � r   d e t . U V i l l   d u   l � g g a   t i l l   a p p l i k a t i o n e n s   s � k v � g   ' % s '   t i l l   m i l j � v a r i a b e l n s   s � k v � g   ( % % P A T H % % ) ? �E d i t o r n   ( a p p l i k a t i o n )   s o m   s t a r t a d e s   f � r   a t t   � p p n a   f i l   ' % s '   a v s l u t a d e s   f � r   t i d i g t .   O m   d e n   i n t e   a v s l u t a d e s   a v   e r ,   k a n   d e t   b e r o   p �   a t t   d e n   e x t e r n a   e d i t o r   � p p n a r   f l e r a   f i l e r   i   e t t   f � n s t e r   ( p r o c e s s ) .   Y t t e r l i g a r e   s t a r t a d e   i n s t a n s e r   a v   e d i t o r n   s k i c k a r   s e d a n   d e n   n y a   f i l e n   t i l l   b e f i n t l i g a   i n s t a n s e r   a v   e d i t o r n   o c h   a v s l u t a r   s i g   o m e d e l b a r t .   F � r   a t t   s t � d j a   d e n n a   t y p   a v   e d i t o r s ,   m � s t e   W i n S C P   a n p a s s a   s i t t   b e t e e n d e ,   i n t e   t a   b o r t   t e m p o r � r   f i l   n � r   p r o c e s s e n   a v s l u t a r ,   u t a n   a t t   b e h � l l a   d e n   s �   l � n g e   W i n S C P   � r   i g � n g .   B e t e e n d e t   k a n   s t � n g a s   a v   g e n o m   a t t   � n d r a   i n s t � l l n i n g a r   f � r   e d i t o r n   ' E x t e r n   e d i t o r   � p p n a r   v a r j e   f i l   i   e t t   s e p a r a t   f � n s t e r   ( p r o c e s s ) ' .   O m   d i n   e d i t o r   i n t e   � r   a v   d e t   h � r   s l a g e t ,   b o r t s e   f r � n   d e t t a   m e d d e l a n d e   o c h   l � t   f i l e n   t a s   b o r t   f r � n   d e n   t e m p o r � r a   k a t a l o g e n   n u . 
   
 V i l l   n i   t a   b o r t   d e n   � p p n a d e   f i l e n   n u ?   ( G e n o m   a t t   t r y c k a   p �   ' N e j '   k o m m e r   d u   a t t   m � j l i g g � r a   d e t   s � r s k i l d a   b e t e e n d e t   o c h   b e h � l l a   f i l e n   i   t e m p o r � r a   m a p p e n . )   � D u   h a r   � s i d o s a t t   f � r v a l d   r i k t n i n g   p �   s y n k r o n i s e r i n g .   S o m   s t a n d a r d   b e s t � m s   r i k t n i n g e n   f r � n   d e n   f i l p a n e l   s o m   v a r   a k t i v   f � r e   k � r n i n g   a v   s y n k r o n i s e r i n g . 
   
 V i l l   d u   a t t   r i k t n i n g e n   d u   v a l d e   s k a   s � t t a s   t i l l   s t a n d a r d ? � V i l l   d u   u t f � r a   f u l l   s y n k r o n i s e r i n g   p �   f j � r r k a t a l o g e n   f � r s t ? 
   
 F u n k t i o n e n   ' H � l l   f j � r r k a t a l o g e n   u p p d a t e r a d '   f u n g e r a r   e n d a s t   k o r r e k t ,   o m   f j � r r k a t a l o g e n   � r   s y n k r o n i s e r a d   m e d   l o k a l   k a t a l o g   i n n a n   d e n   s t a r t a r . 
 1 S � k e r   p �   a t t   d u   v i l l   t a   b o r t   s p a r a d   s e s s i o n   ' % s ' ? � F l e r   � n   % d   k a t a l o g e r   o c h   u n d e r k a t a l o g e r   h i t t a d e s .   B e v a k n i n g   a v   � n d r i n g a r   i   m � n g a   k a t a l o g e r   k a n   s i g n i f i k a n t   m i n s k a   p r e s t a n d a n   p �   d a t o r n . 
   
 V i l l   d u   s k a n n a   f l e r   k a t a l o g e r ,   u p p   t i l l   % d   k a t a l o g e r ? 	 % s   ( % d   s ) 8 S � k e r   p �   a t t   d u   v i l l   f l y t t a   f i l   ' % s '   t i l l   p a p p e r s k o r g e n ? > S � k e r   p �   a t t   d u   v i l l   f l y t t a   % d   v a l d a   f i l e r   t i l l   p a p p e r s k o r g e n ? I F i l e n   h a r   � n d r a t s .   � n d r i n g a r   v i l l   f � r l o r a s ,   o m   f i l e n   l a d d a s   o m .   F o r t s � t t ?  K & o n f i g u r e r a . . . a K a n   i n t e   � p p n a   m o t s v a r a n d e   k a t a l o g   p �   d e n   m o t s a t t a   p a n e l e n . 
   
 V i l l   d u   f � r s � k a   s k a p a   k a t a l o g   ' % s ' ?  L � g g   t i l l   & d e l a d e   b o k m � r k e n �V i l l   d u   s k i c k a   m e d d e l a n d e t   t i l l   W i n S C P : s   w e b b p l a t s ? 
 
 D e t   f i n n s   i n g e n   h j � l p s i d a   a s s o c i e r a d   m e d   m e d d e l a n d e t .   W i n S C P   k a n   s � k a   e f t e r   m e d d e l a n d e t e x t e n   i   d o k u m e n t a t i o n   p �   w e b b p l a t s e n   � t   d i g . 
 
 N o t :   W i n S C P   k o m m e r   a t t   s k i c k a   m e d d e l a n d e t   � v e r   e n   o s � k e r   i n t e r n e t a n s l u t n i n g .   K o n t r o l l e r a   a t t   m e d d e l a n d e t   i n t e   i n n e h � l l e r   n � g o n   i n f o r m a t i o n   s o m   d u   v i l l   s k y d d a ,   s � s o m   n a m n   p �   f i l e r ,   k o n t o n   o c h   v � r d a r . >D i t t   l � s e n o r d   � r   f � r   e n k e l t   o c h   g e r   k a n s k e   i n t e   t i l l r � c k l i g t   m e d   s k y d d   m o t   l e x i k o n   e l l e r   b r u t e - f o r c e   a t t a c k e r . 
   � r   d u   s � k e r   p �   a t t   d u   v i l l   a n v � n d a   d e t ? 
 
 N o t e r a :   b r a   l � s e n o r d   b � r   i n n e h � l l a   m i n s t   s e x   t e c k e n   o c h   b � d e   s t o r a   o c h   s m �   b o k s t � v e r ,   s i f f r o r   o c h   s p e c i a l t e c k e n ,   s o m   a v g r � n s a r e ,   s y m b o l e r ,   b o k s t � v e r   m e d   a c c e n t ,   e t c .                                  W I N _ I N F O R M A T I O N  % s   -   % s  I n g a   s k i l l n a d e r   h i t t a d e s .  � p p n a r   s e s s i o n   ' % s ' 
 % s ' V � n t a r   p �   a t t   d o k u m e n t e t   s k a   s t � n g a s . . . ! % s   ( l a d d a   u p p   m e d   S F T P   e l l e r   S C P ) ! % s   ( l a d d a   u p p   m e d   S F T P   e l l e r   S C P )  L o k a l :   % s 
 F j � r r :   % s    & T o u c h  & K � r     1 % d   f e l   u p p s t o d   v i d   s e n a s t e   o p e r a t i o n e n .   V i s a   d e m ?  F e l   % d   a v   % d : 
 % s  D u   h a r   d e n   s e n a s t e   v e r s i o n e n .  N y   v e r s i o n   % s   h a r   s l � p p t s . % s ! ' % s '   v � r d e   p �   k o m m a n d o & p a r a m e t e r :  ' % s '   k o m m a n d o p a r a m e t e r                        U R L :   P r o t o k o l l e t   % s  A n s l u t e r . . .  F r � g a  F e l  P r o m p t 	 V � n t a r . . .  T a & r / G Z i p . . .  & A r k i v n a m n :  & U n T a r / G Z i p . . .  P a c k a   & u p p   t i l l   k a t a l o g :  & J � m f � r   f i l e r  & G r e p . . .    & S � k   e f t e r   m � n s t e r :  % d   L � s e r   k a t a l o g  B e r � k n a r . . .  
   
 % s 
 L a d d a   & n e r  & K o n t r o l l a   i g e n ; F � r i n s t � l l d   � v e r f � r i n g s i n s t � l l n i n g   ' % s '   v a l d e s   a u t o m a t i s k t . 4 � t e r g �   t i l l   f � r i n s t � l l d   � v e r f � r i n g s i n s t � l l n i n g   ' % s ' . + � t e r g �   t i l l   s t a n d a r d � v e r f � r i n g s i n s t � l l n i n g .  R e g e l   f � r   a u t o m a t i s k t   v a l : 
 % s  & D i s k u t r y m m e s a n v � n d n i n g  A d   H o c  P a u s a  & I n t e r n   e d i t o r �A p p l i k a t i o n   s t a r t a d   f � r   a t t   � p p n a   f i l   ' % s '   s t � n g d e s   f � r   t i d i g t .   O m   d e n   i n t e   s t � n g d e s   a v   d i g ,   d e   k a n   b e r o   p �   a t t   a p p l i k a t i o n e n   � p p n a r   f l e r a   f i l e r   i   e t t   f � n s t e r   ( p r o c e s s ) .   Y t t e r l i g g a r e   s t a r t a d e   i n s t a n s e r   a v   a p p l i k a t i o n e n   s k i c k a r   d �   d e n   n y a   f i l e n   t i l l   b e f i n t l i g   a p p l i k a t i o n   o c h   s t � n g s   o m e d e l b a r t .   W i n S C P   k a n   s t � d j a   s � d a n a   a p p l i k a t i o n e r   e n d a s t   s o m   e x t e r n   e d i t o r . 
   
 O m   d u   v i l l   a n v � n d a   a p p l i k a t i o n e n   f � r   a t t   � p p n a   f i l e r   f r � n   W i n S C P ,   � v e r v � g a   a t t   k o n f i g u r e r a   d e n   s o m   e n   e x t e r n   e d i t o r . 8 R e d i g e r a   ( i n t e r n ) | R e d i g e r a   v a l d a   f i l e r   m e d   i n t e r n   e d i t o r = R e d i g e r a   ( e x t e r n ) | R e d i g e r a   v a l d a   f i l e r   m e d   e x t e r n   e d i t o r   ' % s ' n*   m a t c h a r   e t t   v a l f r i t t   a n t a l   t e c k e n . 
 ?   m a t c h a r   e x a k t   e t t   t e c k e n . 
 [ a b c ]   m a t c h a r   e t t   t e c k e n   f r � n   g r u p p e n . 
 [ a - z ]   m a t c h a r   e t t   t e c k e n   f r � n   i n t e r v a l l e t . 
 > s i z e   m a t c h a r   f i l   s o m   � r   s t � r r e   � n   s t o r l e k e n 
 < s i z e   m a t c h a r   f i l   s o m   � r   m i n d r e   � n   s t o r l e k e n 
 M a s k e r   � r   � t s k i l d a   m e d   s e m i k o l o n   e l l e r   k o m m a t e c k e n . 
 P l a c e r a   e x k l u d e r a d e   m a s k e r   e f t e r   p i p e . 
 E x e m p e l :   * . h t m l ;   p h o t o ? ? . p n g ;   * . z i p > 1 G � M a s k   k a n   f � r l � n g a s   m e d   s � k v � g s m a s k . 
 E x e m p e l :   * / p u b l i c _ h t m l / * . h t m l 
 M a s k   s o m   s l u t a r   m e d   s n e d s t r e c k   m a t c h a r   e n d a s t   k a t a l o g e r . 
 F � r   a t t   m a t c h a   a l l a   k a t a l o g e r   a n v � n d   * / �M � n s t e r : 
 ! !   u t � k a s   t i l l   u t r o p s t e c k e n 
 !   u t � k a s   t i l l   f i l n a m n 
 ! &   u t � k a s   t i l l   l i s t a   m e d   v a l d a   f i l e r   ( c i t a t ,   s p a c e - a v g r � n s a t ) 
 ! /   u t � k a s   t i l l   a k t u e l l   f j � r r s � k v � g 
 ! @   u t � k a s   t i l l   a k t u e l l   s e s s i o n s v � r d n a m n 
 ! U   u t � k a s   t i l l   a k t u e l l   s e s s i o n a s a n v � n d a r n a m n 
 ! P   u t � k a s   t i l l   a k t u e l l   s e s s i o n s l � s e n o r d 
 ! ? p r o m p t [ \ ] ? s t a n d a r d !   u t � k a s   t i l l   a n v � n d a r d e f i n i e r a t   v � r d e   m e d   g i v e n   p r o m p t   o c h   s t a n d a r d   ( a l t e r n a t i v   \   u n d v i k e r   e s c a p i n g ) 
   
 L o k a l t   m � n s t e r k o m m a n d o : 
 ! ^ !   u t � k a s   t i l l   f i l n a m n   f r � n   l o k a l   p a n e l 
   
 E x e m p e l : 
 g r e p   " ! ? M � n s t e r : ? ! "   ! & A A l l a   � v e r f � r i n g a r   i   b a k g r u n d e n   s l u t f � r d e s .   A n s l u t n i n g   a v s l u t a d e s .   L � s n i n g   a v   f j � r r k a t a l o g   a v b r � t s . ( S y n k r o n i s e r a d   b l � d d r i n g   s a t t e s   % s . | p � | a v ' V i s n i n g   a v   d o l d a   f i l e r   s a t t e s   % s . | p � | a v G A u t o m a t i s k   u p p d a t e r i n g   a v   f j � r r k a t a l o g   e f t e r   o p e r a t i o n   s a t t e s   % s . | p � | a v 1 � v e r f � r i n g   i   b a k g r u n d e n   k r � v e r   d i n   u p p m � r k s a m h e t .  � v e r f � r i n g s k �   � r   t o m . M ! Y   � r 
 ! M   m � n a d 
 ! D   d a g 
 ! T   t i d 
 ! @   v � r d n a m n 
 ! S   s e s s i o n s n a m n 
 E x e m p e l :   C : \ ! S ! T . l o g K P a s s i v t   l � g e   m � s t e   v a r a   a k t i v e r a d   n � r   F T P   a n s l u t n i n g   g e n o m   p r o x y   h a r   v a l t s . L U p p d a t e r i n g s k o n t r o l l   f � r   a p p l i k a t i o n e n   � r   t e m p o r � r t   a v s t � n g d .   F � r s � k   s e n a r e .  & G �   t i l l  V a d   � r   n y t t    O p e r a t i o n e n   s l u t f � r d e s  & P r i n t  & A s s o c i e r a d   a p p l i k a t i o n  P �  A v  A u t o P H u v u d l � s e n o r d e t   h a   s a t t s .   D i n a   s p a r a d e   l � s e n o r d   � r   s � k r a d e   g e n o m   A E S   k r y p t e r i n g .  H u v u d l � s e n o r d e t   h a r   � n d r a t s . P D u   h a r   t a g i t   b o r t   d i t t   h u v u d l � s e n o r d .   D i n a   s p a r a d e   l � s e n o r d   s k y d d a s   i n t e   l � n g r e .  H u v u d l � s e n o r d :              W I N _ F O R M S _ S T R I N G S  I n g e n   s e s s i o n s l o g g .  L o g g n i n g   t i l l   f i l   � r   a v s t � n g d . 
 I n g e n   l o g g  S e s s i o n   ' % s '   l o g g  % s   f i l   ' % s '   t i l l   % s :  % s   % d   f i l e r   t i l l   % s :  K o p i e r a  F l y t t a  l o k a l   k a t a l o g  f j � r r k a t a l o g  K o p i e r a  F l y t t a 	 s l � p p   m � l  K o p i e r a  F l y t t a  K o p i e r a r  F l y t t a r  T a r   b o r t  S t � l l e r   i n   i n s t � l l n i n g a r  T e m p o r � r   k a t a l o g  N y   m a p p     	 A v m a r k e r a  M a r k e r a  % d   f i l  % d   f i l e r  % d   m a p p 	 % d   m a p p a r  % d   s y m b o l i s k   l � n k  % d   s y m b o l i s k a   l � n k a r    % s   E g e n s k a p e r  % s ,   . . .   E g e n s k a p e r  A n g e   g i l t i g t   g r u p p n a m n .  A n g e   g i l t i g t   � g a r n a m n .  T i l l b a k a   t i l l   % s  F r a m � t   t i l l   % s      A n s l u t n i n g s t i d  K o m p r i m e r i n g   ( % s )      I n f o r m a t i o n   o m   v a l d   f i l 7 K o m p r i m e r i n g   ( k l i e n t   �   s e r v e r :   % s ,   s e r v e r   �   k l i e n t :   % s )   P � p p n a   s p a r a d   s e s s i o n   ' % s '   ( h � l l   n e r e   S H I F T   f � r   a t t   � p p n a   s e s s i o n   i   n y t t   f � n s t e r )      L i c e n s   f � r   % s                � p p n a   k a t a l o g  H a n t e r a   b o k m � r k e n             
 R a d :   % d / % d 
 K o l u m n :   % d  T e c k e n :   % d   ( 0 x % . 2 x )  � n d r a d  K a n   i n t e   h i t t a   s t r � n g e n   ' % s ' .  T o t a l t   a n t a l   e r s � t t n i n g a r :   % d  G �   t i l l   r a d 
 R a d n u m m e r :  O g i l t i g t   r a d n u m m e r .  R e d i g e r a   l � n k / g e n v � g  L � g g   t i l l   l � n k / g e n v � g  F r � n k o p p l a d .  A n s l u t e r . . .  V � l j   s e s s i o n   ' % s '  L � g g   t i l l   p l a t s p r o f i l  P l a t s p r o f i l n a m n :    F l y t t a   p l a t s p r o f i l  N y t t   m a p p n a m n :  S p a r a   s e s s i o n   s o m  & S p a r a   s e s s i o n   s o m : $ S p a r a   & l � s e n o r d   ( r e k o m m e n d e r a s   i n t e )    K � r   e g e t   k o m m a n d o  K � r   e g e t   k o m m a n d o   ' % s '          K  R 5 % s ,   % d   p t 
 T h e   Q u i c k   B r o w n   F o x   J u m p s   O v e r   T h e   L a z y   D o g  O k � n d    B e r � k n a   k a t a l o g s t o r l e k        A l l m � n n a   i n s t � l l n i n g a r  L a g r a d e   s e s s i o n e r  C a c h a d e   v � r d n y c k l a r  K o n f i g u r a t i o n e n s   I N I - f i l  F i l   m e d   s l u m p f r �  V � l j   l o k a l   k a t a l o g .  F l y t t a r      F l y t t a  H � l l   f j � r r k a t a l o g e n   u p p d a t e r a d % B e h � l l e r   f j � r r k a t a l o g e n   u p p d a t e r a d . . .    T e m p o r � r a   m a p p a r  N y   f i l  R e d i g e r a   f i l  & S k r i v   f i l n a m n : ( D u p l i c a t e   f i l e   ' % s '   t o   r e m o t e   d i r e c t o r y : ' D u p l i c a t e   % d   f i l e s   t o   r e m o t e   d i r e c t o r y :  D u b b l e r a  K o p i e r a r  L � g g   t i l l   e g e t   k o m m a n d o  R e d i g e r a   e g e t   k o m m a n d o  L  F            H � & m t a   f l e r . . .  V � l j   e d i t o r a p p l i k a t i o n . 0 K � r b a r a   f i l e r   ( * . e x e ) | * . e x e | A l l a   f i l e r   ( * . * ) | * . *  % s   a v   % s   i   % s   a v   % s , L � g g   t i l l   f � r i n s t � l l d   � v e r f � r i n g s i n s t � l l n i n g + R e d i g e r a   f � r i n s t � l l d   � v e r f � r i n g s i n s t � l l n i n g 	 S & t a n d a r d  & K o n f i g u r e r a . . .  E g & e t . . .  E g e t   k o m m a n d o  L � g g   t i l l   e d i t o r  R e d i g e r a   e d i t o r  % s ,   B a s e r a s   p �   % s   v e r s i o n   % s  & � p p n a  & K o p i e r a  E n d a s t   & s a m m a   s t o r l e k   N u m b e r   o f   L i c e n s e s :   % s | U n l i m i t e d  P r o d u c t   I D :   % s  % s   ( E x p i r a t i o n   o n   % s )  % s       E d u c a t i o n a l   L i c e n s e  H � m t a r   e g e n s k a p e r    S S H   i m p l e m e n t a t i o n  K r y p t e r i n g s a l g o r i t m  K o m p r i m e r i n g  F i l � v e r f � r i n g s p r o t o k o l l  K a n   � n d r a   r � t t i g h e t e r  K a n   � n d r a   � g a r e / g r u p p  K a n   k � r a   g o d t y c k l i g t   k o m m a n d o " K a n   s k a p a   s y m b o l i s k   l � n k / h � r d   l � n k  K a n   s l �   u p p   a n v � n d a r g r u p p e r  K a n   d u b b l e r a   f j � r r f i l e r   $ � v e r f � r i n g s l � g e   f � r   r e n   t e x t   ( A S C I I ) $ K a n   k o n t r o l l e r a   t i l l g � n g l i g t   u t r y m m e  T o t a l t   a n t a l   b y t e s   p �   e n h e t  L e d i g t   a n t a l   b y t e s   p �   e n h e t   T o t a l t   a n t a l   b y t e s   f � r   a n v � n d a r e  L e d i g a   b y t e s   f � r   a n v � n d a r e  B y t e s   p e r   a l l o k e r i n g s e n h e t  O k � n d  H i t t a   P u T T Y s   p r o g r a m f i l W P u T T Y - p r o g r a m f i l   ( p u t t y . e x e ) | p u t t y . e x e | K � r b a r a   f i l e r   ( * . e x e ) | * . e x e | A l l a   f i l e r   ( * . * ) | * . *  % s   a v   % s | N / A  J � m f � r  S y n k r o n i s e r i n g  A u t e n t i s e r i n g s b a n e r * I N I - f i l   ( * . i n i ) | * . i n i | A l l a   f i l e r   ( * . * ) | * . * ) V � l j   f i l   a t t   e x p o r t e r a   i n s t � l l n i n g a r   t i l l    S & e n s a s t e :   % s 	 S & e n s a s t e  B e r � k n a r   f i l k o n t r o l l s u m m a  K a n   b e r � k n a   f i l k o n t r o l l s u m m a  O k � n d  P r o t o k o l l   s o m   a n v � n d s    O s � k e r   a n s l u t n i n g  S � k e r   a n s l u t n i n g   ( % s )  E n d a s t   p r o t o k o l l k o m m a n d o n  F j � r r s y s t e m  S e s s i o n s p r o t o k o l l      M i n a   d o k u m e n t 	 S k r i v b o r d  K o m m a n d o  S � t t   t i l l   s & t a n d a r d  - -   v a r n a   e f t e r   d e t t a   - -  3 D E S  B l o w f i s h  A E S   ( e n d a s t   S S H - 2 )  D E S  A r c f o u r   ( e n d a s t   S S H - 2 )  - -   v a r n a   e f t e r   d e t t a   - -  D i f f i e - H e l l m a n   g r u p p   1  D i f f i e - H e l l m a n   g r u p p   1 4  D i f f i e - H e l l m a n   g r u p p   u t b y t e  R S A - b a s e r a t   n y c k e l u t b y t e      V � l j   l o k a l   p r o x y a p p l i k a t i o n   � M � n s t e r : 
 \ n   f � r   n y   r a d 
 \ r   f � r   v a g n r e t u r 
 \ t   f � r   t a b 
 \ x X X   f � r   h e x a d e c i m a l   a s c i i k o d 
 \ \   f � r   b a c k s l a s h 
 % v � r d   u t � k a s   t i l l   v � r d n a m n 
 % p o r t   u t � k a s   t i l l   p o r t n u m m e r 
 % u a n v � n d a r e   u t � k a s   t i l l   p r o x y a n v � n d a r n a m n 
 % l � s e n   u t � k a s   t i l l   p r o x y l � s e n o r d 
 % %   f � r   p r o c e n t t e c k e n * S e s s i o n s k a t a l o g   m e d   n a m n   ' % s '   f i n n s   r e d a n . E � r   d u   s � k e r   a t t   d u   v i l l   r a d e r a   s e s s i o n s k a t a l o g   ' % s '   m e d   % d   s e s s i o n e r ? $ K a n   i n t e   r a d e r a   s p e c i a l s e s s i o n   ' % s ' .  S k a p a   s e s s i o n s k a t a l o g  N y t t   m a p p n a m n :   � p p n a   s p a r a d   s e s s i o n k a t a l o g   ' % s '  H o w   t o   p u r c h a s e   a   l i c e n s e . . .  M � l & k a t a l o g : � V i l l   d u   � p p n a   e n   s e p a r a t   s k a l s e s s i o n   f � r   a t t   d u b b l a   f i l e r n a ? 
   
 A k t u e l l   s e s s i o n   s t � d e r   i n t e   d i r e k t   d u b b l i n g   a v   f j � r r f i l e r .   S k i l d a   s k a l s e s s i o n e r   k a n   � p p n a s   f � r   a t t   b e h a n d l a   d u b b l i n g e n .   A l t e r n a t i v t   k a n   d u   d u b b l e r a   f i l e r n a   v i a   l o k a l   t e m p o r � r   k o p i e r i n g .  E d i t o r  % s   ( % s )  % d   d o l d  % d   f i l t r e r a s  F i l t e r � A k t u e l l   s e s s i o n   t i l l � t e r   e n d a s t   f � r � n d r i n g   a v   U I D   � g a n d e t .   D e t   v a r   i n t e   m � j l i g t   a t t   l � s a   U I D   f r � n   k o n t o n a m n e t   " % s " .   S p e c i f i c e r a   U I D   e x p l i c i t   i s t � l l e t .    � v e r f � r   i   & b a k g r u n d e n  % s   ( l � g g   t i l l   i   � v e r f � r i n g s k � )  I n g e n  V � l j   k o r t k o m m a n d o  K o r & t k o m m a n d o : 
 O b e g r � n s a t  H u v u d l � s e n o r d  & N u v a r a n d e   h u v u d l � s e n o r d :  N & y t t   h u v u d l � s e n o r d :  U p p r e p a   h u v u d l � s e n o r d : - S p a r a   & l � s e n o r d   ( s k y d d a s   g e n o m   h u v u d l � s e n o r d ) 	 L e t a   i   % s  S � k 	 S � k e r   . . .  K l a r . 	 A v b r u t e n .    & S t a r t  & S t o p p                                                      W I N _ V A R I A B L E $ C o p y r i g h t   �   2 0 0 0 - 2 0 0 9   M a r t i n   P r i k r y l  h t t p : / / w i n s c p . n e t / " h t t p : / / w i n s c p . n e t / e n g / d o c s / h i s t o r y ' h t t p : / / w i n s c p . n e t / e n g / d o c s / r e q u i r e m e n t s  h t t p : / / w i n s c p . n e t / f o r u m /  h t t p : / / w i n s c p . n e t / u p d a t e s . p h p " h t t p : / / w i n s c p . n e t / e n g / d o w n l o a d . p h p   h t t p : / / w i n s c p . n e t / e n g / d o n a t e . p h p " h t t p : / / w i n s c p . n e t / e n g / d o c s / ? v e r = % s $ h t t p : / / w i n s c p . n e t / e n g / d o c s / % s ? v e r = % s & h t t p : / / w i n s c p . n e t / e n g / t r a n s l a t i o n s . p h p 1 h t t p : / / w i n s c p . n e t / e n g / d o c s / s e a r c h . p h p ? q = % s & v e r = % s                  A n s l u t e n 0 A n s l u t e n   m e d   % s .   V � n t a r   p �   v � l k o m s t m e d d e l a n d e . . .   * A n s l u t e n   m e d   % s ,   f � r m e d l a r   S S L - k o p p l i n g . . .  A n s l u t e r   t i l l   % s   . . .  L i s t i n g   a v   k a t a l o g e r   l y c k a d  K o p p l a r   i f r � n   s e r v e r    s t a r t a r   n e r l a d d n i n g   a v   % s  N e r l a d d n i n g   l y c k a d   * F � r s � k e r   a t t   a n s l u t a   % s   g e n o m   F T P   p r o x y . . .              � t e r f � r   l i s t i n g   a v   k a t a l o g e r . . . 7 S S L - k o p p l i n g   u p p r � t t a d .   V � n t a r   p �   v � l k o m s t m e d d e l a n d e . . .  S S L - k o p p l i n g   u p p r � t t a d  S t a r t a r   u p p l a d d n i n g   a v   % s  U p p l a d d n i n g   l y c k a d                               5 K u n d e   i n t e   s k a p a   s o c k e t   i   d e n   a n g i v n a   p o r t i n t e r v a l l e t    K a n   i n t e   u p p r � t t a   S S L - k o p p l i n g   & K u n d e   i n t e   � t e r f �   l i s t i n g   a v   k a t a l o g e r     # K a n   i n t e   i n i t i a l i s e r a   S S L - b i b l i o t e k       , � v e r f � r i n g s t u n n e l   k a n   i n t e   � p p n a s .   O r s a k :   % s    K a n   i n t e   a v g � r a   v � r d n a m n > � t e r u p p t a g n i n g s k o m m a n d o   s t � d s   i n t e   a v   s e r v e r ,   s k r i v a   � v e r   f i l . I P a u s k o m m a n d o   s t � d s   i n t e   a v   s e r v e r ,   m e n   l o k a l   o c h   f j � r r f i l s t o r l e k   � r   l i k a . , O f � r m � g e n   a t t   s k i c k a   k o m m a n d o .   K o p p l a   i f r � n .    P e e r   c e r t i f i k a t   f � r k a s t a s    N e r l a d d n i n g   a v b r u t e n                      F i l e n   f i n n s   r e d a n          P r o x y   k r � v e r   a u t e n t i s e r i n g P N � d v � n d i g   a u t e n t i s e r i n g s t y p   r a p p o r t e r a d   a v   p r o x y s e r v e r   � r   o k � n d   e l l e r   s t � d s   i n t e % K a n   i n t e   a v g � r a   v � r d   t i l l   p r o x y s e r v e r ! K a n   i n t e   a n s l u t a   t i l l   p r o x y s e r v e r C B e g � r a n   f r � n   p r o x y   m i s s l y c k a d e s ,   k a n   i n t e   a n s l u t a   g e n o m   p r o x y s e r v e r                        T i m o u t   d e t e k t e r a d .  U p p l a d d n i n g   a v b r u t e n            K u n d e   i n t e   s � t t a   f i l p e k a r e  O k � n t   f e l   i   S S L - l a g r e t % K u n d e   i n t e   v e r i f i e r a   S S L - c e r t i f i k a t e t                                               , � v e r s � t t n i n g :   A .   P e t t e r s s o n   < a z @ k t h . s e >   2 0 0 8                          a n   u n n a m e d   f i l e                      N o   e r r o r   m e s s a g e   i s   a v a i l a b l e . ' A n   u n s u p p o r t e d   o p e r a t i o n   w a s   a t t e m p t e d . $ A   r e q u i r e d   r e s o u r c e   w a s   u n a v a i l a b l e .  O u t   o f   m e m o r y .  A n   u n k n o w n   e r r o r   h a s   o c c u r r e d .                                        F a i l e d   t o   l a u n c h   h e l p .  I n t e r n a l   a p p l i c a t i o n   e r r o r .  C o m m a n d   f a i l e d . ) I n s u f f i c i e n t   m e m o r y   t o   p e r f o r m   o p e r a t i o n . P S y s t e m   r e g i s t r y   e n t r i e s   h a v e   b e e n   r e m o v e d   a n d   t h e   I N I   f i l e   ( i f   a n y )   w a s   d e l e t e d . B N o t   a l l   o f   t h e   s y s t e m   r e g i s t r y   e n t r i e s   ( o r   I N I   f i l e )   w e r e   r e m o v e d . F T h i s   p r o g r a m   r e q u i r e s   t h e   f i l e   % s ,   w h i c h   w a s   n o t   f o u n d   o n   t h i s   s y s t e m . t T h i s   p r o g r a m   i s   l i n k e d   t o   t h e   m i s s i n g   e x p o r t   % s   i n   t h e   f i l e   % s .   T h i s   m a c h i n e   m a y   h a v e   a n   i n c o m p a t i b l e   v e r s i o n   o f   % s .      P l e a s e   e n t e r   a n   i n t e g e r .  P l e a s e   e n t e r   a   n u m b e r . * P l e a s e   e n t e r   a n   i n t e g e r   b e t w e e n   % 1   a n d   % 2 . ( P l e a s e   e n t e r   a   n u m b e r   b e t w e e n   % 1   a n d   % 2 . ( P l e a s e   e n t e r   n o   m o r e   t h a n   % 1   c h a r a c t e r s .  P l e a s e   s e l e c t   a   b u t t o n . * P l e a s e   e n t e r   a n   i n t e g e r   b e t w e e n   0   a n d   2 5 5 .   P l e a s e   e n t e r   a   p o s i t i v e   i n t e g e r .   P l e a s e   e n t e r   a   d a t e   a n d / o r   t i m e .  P l e a s e   e n t e r   a   c u r r e n c y .                U n e x p e c t e d   f i l e   f o r m a t . V % 1 
 C a n n o t   f i n d   t h i s   f i l e . 
 P l e a s e   v e r i f y   t h a t   t h e   c o r r e c t   p a t h   a n d   f i l e   n a m e   a r e   g i v e n .  D e s t i n a t i o n   d i s k   d r i v e   i s   f u l l . 5 U n a b l e   t o   r e a d   f r o m   % 1 ,   i t   i s   o p e n e d   b y   s o m e o n e   e l s e . A U n a b l e   t o   w r i t e   t o   % 1 ,   i t   i s   r e a d - o n l y   o r   o p e n e d   b y   s o m e o n e   e l s e . . A n   u n e x p e c t e d   e r r o r   o c c u r r e d   w h i l e   r e a d i n g   % 1 . . A n   u n e x p e c t e d   e r r o r   o c c u r r e d   w h i l e   w r i t i n g   % 1 .                                           # U n a b l e   t o   r e a d   w r i t e - o n l y   p r o p e r t y . # U n a b l e   t o   w r i t e   r e a d - o n l y   p r o p e r t y .      N o   e r r o r   o c c u r r e d . - A n   u n k n o w n   e r r o r   o c c u r r e d   w h i l e   a c c e s s i n g   % 1 .  % 1   w a s   n o t   f o u n d .  % 1   c o n t a i n s   a n   i n v a l i d   p a t h . = % 1   c o u l d   n o t   b e   o p e n e d   b e c a u s e   t h e r e   a r e   t o o   m a n y   o p e n   f i l e s .  A c c e s s   t o   % 1   w a s   d e n i e d . . A n   i n v a l i d   f i l e   h a n d l e   w a s   a s s o c i a t e d   w i t h   % 1 . < % 1   c o u l d   n o t   b e   r e m o v e d   b e c a u s e   i t   i s   t h e   c u r r e n t   d i r e c t o r y . 6 % 1   c o u l d   n o t   b e   c r e a t e d   b e c a u s e   t h e   d i r e c t o r y   i s   f u l l .  S e e k   f a i l e d   o n   % 1 5 A   h a r d w a r e   I / O   e r r o r   w a s   r e p o r t e d   w h i l e   a c c e s s i n g   % 1 . 0 A   s h a r i n g   v i o l a t i o n   o c c u r r e d   w h i l e   a c c e s s i n g   % 1 . 0 A   l o c k i n g   v i o l a t i o n   o c c u r r e d   w h i l e   a c c e s s i n g   % 1 .  D i s k   f u l l   w h i l e   a c c e s s i n g   % 1 . . A n   a t t e m p t   w a s   m a d e   t o   a c c e s s   % 1   p a s t   i t s   e n d .    N o   e r r o r   o c c u r r e d . - A n   u n k n o w n   e r r o r   o c c u r r e d   w h i l e   a c c e s s i n g   % 1 . / A n   a t t e m p t   w a s   m a d e   t o   w r i t e   t o   t h e   r e a d i n g   % 1 . . A n   a t t e m p t   w a s   m a d e   t o   a c c e s s   % 1   p a s t   i t s   e n d . 0 A n   a t t e m p t   w a s   m a d e   t o   r e a d   f r o m   t h e   w r i t i n g   % 1 .  % 1   h a s   a   b a d   f o r m a t . " % 1   c o n t a i n e d   a n   u n e x p e c t e d   o b j e c t .   % 1   c o n t a i n s   a n   i n c o r r e c t   s c h e m a .                 / M e n u   ' % s '   i s   a l r e a d y   b e i n g   u s e d   b y   a n o t h e r   f o r m  P i c t u r e :    ( % d x % d )  P r e v i e w  C a n n o t   o p e n   A V I  D o c k e d   c o n t r o l   m u s t   h a v e   a   n a m e % E r r o r   r e m o v i n g   c o n t r o l   f r o m   d o c k   t r e e    -   D o c k   z o n e   n o t   f o u n d    -   D o c k   z o n e   h a s   n o   c o n t r o l , M u l t i s e l e c t   m o d e   m u s t   b e   o n   f o r   t h i s   f e a t u r e 	 S e p a r a t o r  E r r o r   s e t t i n g   % s . C o u n t 8 L i s t b o x   ( % s )   s t y l e   m u s t   b e   v i r t u a l   i n   o r d e r   t o   s e t   C o u n t          R i g h t  D o w n  I n s  D e l  S h i f t +  C t r l +  A l t +  ( N o n e )  V a l u e   m u s t   b e   b e t w e e n   % d   a n d   % d  A l l  U n a b l e   t o   i n s e r t   a   l i n e  I n v a l i d   c l i p b o a r d   f o r m a t   C l i p b o a r d   d o e s   n o t   s u p p o r t   I c o n s  C a n n o t   o p e n   c l i p b o a r d  T e x t   e x c e e d s   m e m o   c a p a c i t y . T h e r e   i s   n o   d e f a u l t   p r i n t e r   c u r r e n t l y   s e l e c t e d  & F � r s � k   i g e n 	 & I g n o r e r a  & A l l a  N & e j   t i l l   a l l a  J & a   t i l l   a l l a  B k S p  T a b  E s c  E n t e r  S p a c e  P g U p  P g D n  E n d  H o m e  L e f t  U p 	 M e t a f i l e s  E n h a n c e d   M e t a f i l e s  I c o n s  B i t m a p s  O g i l t i g t   i n p u t v � r d e 9 O g i l t i g t   i n p u t v � r d e .   A n v � n d   E S C   f � r   a t t   a v b r y t a   � n d r i n g a r  V a r n i n g  F e l  I n f o r m a t i o n  B e k r � f t a  & J a  & N e j  O K  A v b r y t  & H j � l p  & A v b r y t  P r i n t e r   s e l e c t e d   i s   n o t   v a l i d  % s   o n   % s @ G r o u p I n d e x   c a n n o t   b e   l e s s   t h a n   a   p r e v i o u s   m e n u   i t e m ' s   G r o u p I n d e x 5 C a n n o t   c r e a t e   f o r m .   N o   M D I   f o r m s   a r e   c u r r e n t l y   a c t i v e * A   c o n t r o l   c a n n o t   h a v e   i t s e l f   a s   i t s   p a r e n t  O K  A v b r y t  & Y e s  & N o  & H e l p  & C l o s e  & I g n o r e  & R e t r y  A b o r t  & A l l  C a n n o t   d r a g   a   f o r m ( F a i l e d   t o   w r i t e   I m a g e L i s t   d a t a   t o   s t r e a m $ E r r o r   c r e a t i n g   w i n d o w   d e v i c e   c o n t e x t  E r r o r   c r e a t i n g   w i n d o w   c l a s s + C a n n o t   f o c u s   a   d i s a b l e d   o r   i n v i s i b l e   w i n d o w ! C o n t r o l   ' % s '   h a s   n o   p a r e n t   w i n d o w $ P a r e n t   g i v e n   i s   n o t   a   p a r e n t   o f   ' % s '  C a n n o t   h i d e   a n   M D I   C h i l d   F o r m ) C a n n o t   c h a n g e   V i s i b l e   i n   O n S h o w   o r   O n H i d e " C a n n o t   m a k e   a   v i s i b l e   w i n d o w   m o d a l  % s   p r o p e r t y   o u t   o f   r a n g e  M e n u   i n d e x   o u t   o f   r a n g e  M e n u   i n s e r t e d   t w i c e  S u b - m e n u   i s   n o t   i n   m e n u  N o t   e n o u g h   t i m e r s   a v a i l a b l e ! P r i n t e r   i s   n o t   c u r r e n t l y   p r i n t i n g  P r i n t i n g   i n   p r o g r e s s  B i t m a p   i m a g e   i s   n o t   v a l i d  I c o n   i m a g e   i s   n o t   v a l i d  M e t a f i l e   i s   n o t   v a l i d  I n v a l i d   p i x e l   f o r m a t  I n v a l i d   i m a g e  S c a n   l i n e   i n d e x   o u t   o f   r a n g e ! C a n n o t   c h a n g e   t h e   s i z e   o f   a n   i c o n $ U n k n o w n   p i c t u r e   f i l e   e x t e n s i o n   ( . % s )  U n s u p p o r t e d   c l i p b o a r d   f o r m a t  O u t   o f   s y s t e m   r e s o u r c e s  C a n v a s   d o e s   n o t   a l l o w   d r a w i n g  I n v a l i d   i m a g e   s i z e  I n v a l i d   I m a g e L i s t  U n a b l e   t o   R e p l a c e   I m a g e  I n v a l i d   I m a g e L i s t   I n d e x ) F a i l e d   t o   r e a d   I m a g e L i s t   d a t a   f r o m   s t r e a m     F a i l e d   t o   d e l e t e   t a b   a t   i n d e x   % d " F a i l e d   t o   r e t r i e v e   t a b   a t   i n d e x   % d   F a i l e d   t o   g e t   o b j e c t   a t   i n d e x   % d " F a i l e d   t o   s e t   t a b   " % s "   a t   i n d e x   % d   F a i l e d   t o   s e t   o b j e c t   a t   i n d e x   % d < M u l t i L i n e   m u s t   b e   T r u e   w h e n   T a b P o s i t i o n   i s   t p L e f t   o r   t p R i g h t  I n v a l i d   i n d e x  U n a b l e   t o   i n s e r t   a n   i t e m  I n v a l i d   o w n e r  R i c h E d i t   l i n e   i n s e r t i o n   e r r o r  F a i l e d   t o   L o a d   S t r e a m  F a i l e d   t o   S a v e   S t r e a m E % d   i s   a n   i n v a l i d   P a g e I n d e x   v a l u e .     P a g e I n d e x   m u s t   b e   b e t w e e n   0   a n d   % d = T h i s   c o n t r o l   r e q u i r e s   v e r s i o n   4 . 7 0   o r   g r e a t e r   o f   C O M C T L 3 2 . D L L 0 T a b   p o s i t i o n   i n c o m p a t i b l e   w i t h   c u r r e n t   t a b   s t y l e 0 T a b   s t y l e   i n c o m p a t i b l e   w i t h   c u r r e n t   t a b   p o s i t i o n    M o n d a y  T u e s d a y 	 W e d n e s d a y  T h u r s d a y  F r i d a y  S a t u r d a y  U n a b l e   t o   c r e a t e   d i r e c t o r y  T o o l b a r   i t e m   i n d e x   o u t   o f   r a n g e  T o o l b a r   i t e m   a l r e a d y   i n s e r t e d ? A n   i t e m   v i e w e r   a s s o c i a t e d   t h e   s p e c i f i e d   i t e m   c o u l d   n o t   b e   f o u n d  M o r e   B u t t o n s | J A   T T B D o c k   c o n t r o l   c a n n o t   b e   p l a c e d   i n s i d e   a   t o o l   w i n d o w   o r   a n o t h e r   T T B D o c k C C a n n o t   c h a n g e   P o s i t i o n   o f   a   T T B D o c k   i f   i t   a l r e a d y   c o n t a i n s   c o n t r o l s G C a n n o t   s a v e   d o c k a b l e   w i n d o w ' s   p o s i t i o n   b e c a u s e   N a m e   p r o p e r t y   i s   n o t   s e t O C a n n o t   s a v e   d o c k a b l e   w i n d o w ' s   p o s i t i o n   b e c a u s e   D o c k e d T o ' s   N a m e   p r o p e r t y   n o t   s e t  F a i l e d   t o   c l e a r   t a b   c o n t r o l  M a y  J u n e  J u l y  A u g u s t 	 S e p t e m b e r  O c t o b e r  N o v e m b e r  D e c e m b e r  S u n  M o n  T u e  W e d  T h u  F r i  S a t  S u n d a y  J a n  F e b  M a r  A p r  M a y  J u n  J u l  A u g  S e p  O c t  N o v  D e c  J a n u a r y  F e b r u a r y  M a r c h  A p r i l   5 C o u l d   n o t   c o n v e r t   v a r i a n t   o f   t y p e   ( % s )   i n t o   t y p e   ( % s ) = O v e r f l o w   w h i l e   c o n v e r t i n g   v a r i a n t   o f   t y p e   ( % s )   i n t o   t y p e   ( % s )  V a r i a n t   o v e r f l o w  I n v a l i d   a r g u m e n t  I n v a l i d   v a r i a n t   t y p e  O p e r a t i o n   n o t   s u p p o r t e d  U n e x p e c t e d   v a r i a n t   e r r o r  E x t e r n a l   e x c e p t i o n   % x  A s s e r t i o n   f a i l e d  I n t e r f a c e   n o t   s u p p o r t e d  E x c e p t i o n   i n   s a f e c a l l   m e t h o d  % s   ( % s ,   l i n e   % d )  A b s t r a c t   E r r o r ? A c c e s s   v i o l a t i o n   a t   a d d r e s s   % p   i n   m o d u l e   ' % s ' .   % s   o f   a d d r e s s   % p  S y s t e m f e l .     K o d :   % d .  
 % s * E t t   a n r o p   t i l l   e n   O S   f u n k t i o n   m i s s l y c k a d e s ( E x c e p t i o n   % s   i n   m o d u l e   % s   a t   % p .  
 % s % s  
  A p p l i c a t i o n   E r r o r 1 F o r m a t   ' % s '   i n v a l i d   o r   i n c o m p a t i b l e   w i t h   a r g u m e n t  N o   a r g u m e n t   f o r   f o r m a t   ' % s ' " V a r i a n t   m e t h o d   c a l l s   n o t   s u p p o r t e d  R e a d  W r i t e  F o r m a t   s t r i n g   t o o   l o n g  E r r o r   c r e a t i n g   v a r i a n t   a r r a y ! V a r i a n t   a r r a y   i n d e x   o u t   o f   b o u n d s  V a r i a n t   a r r a y   i s   l o c k e d  I n v a l i d   v a r i a n t   t y p e   c o n v e r s i o n  I n v a l i d   v a r i a n t   o p e r a t i o n ! I n v a l i d   v a r i a n t   o p e r a t i o n   ( $ % . 8 x )  V a r i a n t   i s   n o t   a n   a r r a y  I n v a l i d   N U L L   v a r i a n t   o p e r a t i o n 	 D i s k   f u l l  I n v a l i d   n u m e r i c   i n p u t  D i v i s i o n   b y   z e r o  R a n g e   c h e c k   e r r o r  I n t e g e r   o v e r f l o w   I n v a l i d   f l o a t i n g   p o i n t   o p e r a t i o n  F l o a t i n g   p o i n t   d i v i s i o n   b y   z e r o  F l o a t i n g   p o i n t   o v e r f l o w  F l o a t i n g   p o i n t   u n d e r f l o w  I n v a l i d   p o i n t e r   o p e r a t i o n  I n v a l i d   c l a s s   t y p e c a s t 0 A c c e s s   v i o l a t i o n   a t   a d d r e s s   % p .   % s   o f   a d d r e s s   % p  S t a c k   o v e r f l o w  C o n t r o l - C   h i t  P r i v i l e g e d   i n s t r u c t i o n  O p e r a t i o n   a b o r t e d / V a r i a n t   d o e s   n o t   r e f e r e n c e   a n   a u t o m a t i o n   o b j e c t 7 D i s p a t c h   m e t h o d s   d o   n o t   s u p p o r t   m o r e   t h a n   6 4   p a r a m e t e r s ! ' % s '   i s   n o t   a   v a l i d   i n t e g e r   v a l u e ( ' % s '   i s   n o t   a   v a l i d   f l o a t i n g   p o i n t   v a l u e  ' % s '   � r   i n g e t   g i l t i g t   d a t u m  ' % s '   � r   i n g e n   g i l t i g   t i d # ' % s '   � r   i n g e t   g i l t i g t   d a t u m   o c h   t i d  I n v a l i d   a r g u m e n t   t o   t i m e   e n c o d e  I n v a l i d   a r g u m e n t   t o   d a t e   e n c o d e  O u t   o f   m e m o r y  I / O   e r r o r   % d  F i l e   n o t   f o u n d  I n v a l i d   f i l e n a m e  T o o   m a n y   o p e n   f i l e s  F i l e   a c c e s s   d e n i e d  R e a d   b e y o n d   e n d   o f   f i l e  E r r o r   r e a d i n g   % s % s % s :   % s  S t r e a m   r e a d   e r r o r  P r o p e r t y   i s   r e a d - o n l y  F a i l e d   t o   c r e a t e   k e y   % s  F a i l e d   t o   g e t   d a t a   f o r   ' % s '  I n v a l i d   c o m p o n e n t   r e g i s t r a t i o n  F a i l e d   t o   s e t   d a t a   f o r   ' % s '  R e s o u r c e   % s   n o t   f o u n d  % s . S e e k   n o t   i m p l e m e n t e d $ O p e r a t i o n   n o t   a l l o w e d   o n   s o r t e d   l i s t   T o o   m a n y   r o w s   o r   c o l u m n s   d e l e t e d $ % s   n o t   i n   a   c l a s s   r e g i s t r a t i o n   g r o u p  P r o p e r t y   % s   d o e s   n o t   e x i s t  S t r e a m   w r i t e   e r r o r  O L E   e r r o r   % . 8 x . M e t h o d   ' % s '   n o t   s u p p o r t e d   b y   a u t o m a t i o n   o b j e c t   + F i x e d   r o w   c o u n t   m u s t   b e   l e s s   t h a n   r o w   c o u n t  C a n n o t   o p e n   f i l e   % s  G r i d   t o o   l a r g e   f o r   o p e r a t i o n  G r i d   i n d e x   o u t   o f   r a n g e  U n a b l e   t o   w r i t e   t o   % s  I n v a l i d   s t r e a m   f o r m a t  ' % s '   i s   a n   i n v a l i d   m a s k   a t   ( % d ) $ ' ' % s ' '   i s   n o t   a   v a l i d   c o m p o n e n t   n a m e  I n v a l i d   p r o p e r t y   v a l u e  I n v a l i d   p r o p e r t y   p a t h  I n v a l i d   p r o p e r t y   v a l u e  I n v a l i d   d a t a   t y p e   f o r   ' % s '   L i s t   c a p a c i t y   o u t   o f   b o u n d s   ( % d )  L i s t   c o u n t   o u t   o f   b o u n d s   ( % d )  L i s t   i n d e x   o u t   o f   b o u n d s   ( % d ) + O u t   o f   m e m o r y   w h i l e   e x p a n d i n g   m e m o r y   s t r e a m " U n a b l e   t o   f i n d   a   T a b l e   o f   C o n t e n t s  N o   h e l p   f o u n d   f o r   % s # N o   c o n t e x t - s e n s i t i v e   h e l p   i n s t a l l e d $ N o   t o p i c - b a s e d   h e l p   s y s t e m   i n s t a l l e d  A n c e s t o r   f o r   ' % s '   n o t   f o u n d  C a n n o t   a s s i g n   a   % s   t o   a   % s  B i t s   i n d e x   o u t   o f   r a n g e * C a n ' t   w r i t e   t o   a   r e a d - o n l y   r e s o u r c e   s t r e a m E C h e c k S y n c h r o n i z e   c a l l e d   f r o m   t h r e a d   $ % x ,   w h i c h   i s   N O T   t h e   m a i n   t h r e a d  C l a s s   % s   n o t   f o u n d  A   c l a s s   n a m e d   % s   a l r e a d y   e x i s t s % L i s t   d o e s   n o t   a l l o w   d u p l i c a t e s   ( $ 0 % x ) # A   c o m p o n e n t   n a m e d   % s   a l r e a d y   e x i s t s % S t r i n g   l i s t   d o e s   n o t   a l l o w   d u p l i c a t e s  C a n n o t   c r e a t e   f i l e   % s 1 F i x e d   c o l u m n   c o u n t   m u s t   b e   l e s s   t h a n   c o l u m n   c o u n t % F i l n a m n e t   i n n e h � l l e r   o g i l t i g a   t e c k e n :  F i l   % s  % u   F i l e r  % u   K a t a l o g e r  H u v u d k a t a l o g * K a n   i n t e   a v s l u t a   t r � d   f � r   i k o n u p p d a t e r i n g .  D r a S l � p p   f e l :   % d  E n h e t   ' % s : '   � r   i n t e   k l a r .  K a t a l o g e n   ' % s '   f i n n s   i n t e .  /   < r o o t >  R � t t i g h e t e r  � g a r e  G r u p p  M � l   l � n k  F i l t y p  D r a g & d r o p   e r r o r :   % d 	 \ / : * ? " < > |    ' N e w   n a m e   c o n t a i n s   i n v a l i d   c h a r a c t e r s   % s  F i l o p e r a t i o n # K a n   i n t e   h i t t a   n � g o n   g i l t i g   s � k v � g .  U N C   s � k v � g a r   s t � d s   i n t e .  % s   � r   e n   o g i l t i g   e n h e t s b o k s t a v .  N a m n  S t o r l e k  F i l t y p  � n d r a d  A t t r  E x t  K a n   i n t e   � p p n a   f i l :   ) K a n   i n t e   b y t a   n a m n   p �   f i l   e l l e r   k a t a l o g :    F i l e n   f i n n s   r e d a n :      & K o p i e r a   h i t  & F l y t t a   h i t  & S k a p a   g e n v � g   h i t  & A v b r y t  B l � d d r a  A l l a   f i l e r   ( * . * ) | * . *  O g i l t i g t   f i l n a m n   -   % s  S o c k e t   e r r o r   ( % s )  T i m e o u t 	 O k � n t   f e l  R e c e i v e d   r e s p o n s e   % d   % s   f r o m   % s " E x c e e d e d   m a x i m a l   r e d i r e c t   l i m i e   % d  F i l s y s t e m s o p e r a t i o n 	 \ / : * ? " < > |     F i l e s y s t e m   O p e r a t i o n #x]#���C�@&��TPF0TAboutDialogAboutDialogLeftuTop{HelpType	htKeywordHelpKeywordui_aboutBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption	Om WinSCPClientHeight�ClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameMS Sans Serif
Font.Style OldCreateOrder	PositionpoMainFormCenter
DesignSize�� PixelsPerInch`
TextHeight TLabelApplicationLabelLeftHTopWidth4HeightCaptionApplication  TLabelVersionLabelLeftHTopWidth~HeightCaptionVersion 2.0.0 (Build 12) XX  TLabelWinSCPCopyrightLabelLeftHTop8Width� HeightCaption$Copyright � 2000-2003 Martin Prikryl  TLabelProductSpecificMessageLabelLeftHTopdWidthHeightCaption4F�r att skicka in kommentarer och rapportera buggar:  TLabelTranslatorLabelLeftHTop� WidthIHeightCaptionTranslatorLabel  TImageImageLeftTopWidth1Height Center	Picture.Data
� TIcon         h  v        �	  �         �  f  **         00     �%  <  @@     (B  �a  ��     ( �  (                                     jjj�iii�iii�iii�iii�iii�jjj�E�E�T�T�^�_�i�i�s�t�~�~���������k�kXiii���������������������iii�2�4aE�E�����������-�-�����iii���������������������iii��D 2�4aD�E��� �� �� ��������iii���������������������iii��D 0�2;=�>�	�
� �� �� ����~�~�jjj�iii�iii�iii�iii�iii�jjj�� 7)�*��� �� �� �� ����s�t��D fff������D ����fff�]�[��	�� �� �� ��	�
�����i�i��u%	fff������D ����fff�]���� �� �� ����=�>�D�E���^�_��}8�fff�������������fff��z	�/�� �� ��	��(�*�-�.@5�7[E�F�T�T��A��sg�fff�fff�fff�q^��o ��v �-�������<�D �D 5�7[D�E��G��a��}9��5��l��f ��j ��o ��{	�Z��X�^�D �D �D �D 2�3�M��R��X��^	��] ��a ��f ��r����9�D �D �D �D �D �D �R��M��O ��S ��X ��] ��l��*��}!:�D �D �D �D �D �D �D ��X��I��J ��O ��S ��^	��5��}-:�D �D �D �D �D �D �D �D �^��E��E ��J ��O ��X��}9��}2T�D �D �D �D �D �D �D �D �~[��X%��E��I��M��R��a��~:��{0S�D �D �D �D �D �D �D �rOO�~[��^���X��R��M��G��A��}8��u%	�D �D �D �D �D �D       �  �     �   �          ?      �  �  �   �  �  (      0                              ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �Հo�suR�V�M�Q�L�P�L�P�K�P�L�Q�Y�`�'=':   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���b�f��� � � � � � � � � � �� �m�r�   ��� ��� ��� ���                               ^�a��� � � � � � ���>�>�m�r�   ��� ��� ��� ���    CCC"777A111I111I444I444I777J777J777J999LRlTa>�A� � � � ���4�4�>�>�n�q�   ��� ��� ��� ��� ��� ttt�\\\�ggg�fff�mmm�www�zzz�yyy�}}}�����V�X��� � ���*�*�3�3�=�=�m�q�   ��� ��� ��� ��� ���+DDD�(((�222�???�???�===�EEE�CCC�KMK�I}J� �!�������)�)�3�3�<�<�n�q�   ��� ��� ��� ��� ���+JJJ�,,,�777�GGG�HHH�EEE�PPP�MMM�I]I�?u@�6�7�'�(�'�(�!�"�C�D�;�;�<�<�n�q�   ��� ��� ��� ��� ���*GGG�333�>>>�NNN�QQQ�MMM�\\\�VVV�Y]Y�VsW�Q�R�B�C�:�;�L�N�k�nfv�x�D�D�p�s�   
��� ��� ��� ��� ���)AAA�999�DDD�TTT�YYY�SSS�fff�___�ddd�ptp�o�p�Z�[�\�]�����   ���z�}�}び   ��� ��� ��� ��� ���)KKK�@@@�III�ZZZ�```�XXX�ppp�hhh�kkk�}}}�����w�x�x�y�����   ��� ��������� ��� ��� ��� ��� ���(OOO�GGG�MMM�___�ccc�]]]�zzz�qqq�sss�������������xxx�����   ��� ��� ��� ��� ��� ��� ��� ��� ���&PPP�MMM�RRR�bbb�eee�aaa�����xxx�|||���������������������   ��� ��� ��� ���          ��� ���ZZZ�TTT�VVV�eee�ggg�fff�����������������������������v   ��� ��� ��� ��� udW0)$      ������w���򦦦��������Ͷ��������������ƭ������������������"   ��� ��� ��� ��� �uf�f�   �|b��CrwlZ���������GD<Y            	��������eee�      ��� ��� ��� ��� ��� ��R��q��a�r\I:�F��} �|mW���������lX0jRF+   ���    	��������eee�      ��� ��� ��� ��� ��� �L��i ��p��@��v ��x ��mU����������n;��oO         ��������eee�      ��� ��� ��� ��� ��� �G��d ��i ��m ��r ��xËnO���������qj`�   '      /�����ccc�      ��� ��� ��� ��� ��� �C��` ��d ��i ��r��x
��}1թ�����������kkk�jjj�jjj�qqq򨨨�����^^^�   ��� ��� ��� ��� ��� ��� �}>��[ ��` ��j
��q��s
��4؎�������������������������������ggg�      ��� ��� ��� ��� ��� ��� �y;��V ��d��l��m��o
��t��s�zzyā��쒒�򅅅�ttt�lll�eee�+++   ��� ��� ��� ��� ��� ��� ��� ށJr�_��f��h��j��k��m��r��f�(!   	               ��� ��� ��� ��� ��� ��� ��� ��� ��cބN��D���B��B��B��B���C���b�䵔   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �� �� �� �� �  �  �  �  �  �  �  �  � ? � ? �| |  <  <      �  � �� �� (       @                              ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���          
                                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    +t�{Ql�qhg�nme�loc�jqa�gt_�ev\�ct/A   *      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��>h�l�*�,�"�$�"�$�"�$�"�$�"�$�"�%�$�&�Q�V�i�p�   (   ��� ��� ��� ��� ��� ��� ��� ���                               f�fw�|��� � � � � � � � � � � � � � ���m�p�@lFP   ��� ��� ��� ��� ��� ���             	   	   	   	   	   	   	   	   	   	(;(t�y��� � � � � � � � � � ���=�=�I�I�{ނ�   ��� ��� ��� ��� ���             !   %   &   &   &   &   &   &   &   &   &   &+q�t��� � � � � � ���5�5�<�<�D�D�~ᄺ   ��� ��� ��� ��� ���    rrr���^vvv�zzz�vvv�vvv�zzz������������������������������O�Q� � � � � � ���-�-�5�5�<�<�D�D�ⅸ   ��� ��� ��� ��� ���    ���rTTT�FFF�PPP�RRR�PPP�VVV�___�eee�ggg�fff�jjj�ooo�w}w�U�W��� � � � ���&�&�-�-�4�4�<�<�C�C��ᄷ   ��� ��� ��� ��� ���    ����111�&&&�000�666�>>>�===�;;;�???�DDD�BBB�FFF�QUQ�J�K� �!���	�
�	�	���&�&�-�-�4�4�;�;�C�C��ᅶ   ��� ��� ��� ��� ���    ����444�'''�333�:::�FFF�EEE�AAA�FFF�MMM�JJJ�KLK�HkI�6x7�/�0�"�#���!�"���%�%�,�,�4�4�;�;�B�B��↵   ��� ��� ��� ��� ���    ����777�+++�999�>>>�KKK�MMM�GGG�NNN�UUU�PPP�OWO�IfJ�GwH�A�B�5�6�1�2�.�/�)�*�9�9����B�C�;�;�B�B��㈲   ��� ��� ��� ��� ���    ����555�000�@@@�CCC�QQQ�TTT�LLL�SSS�]]]�XXX�YYY�[f[�Zw[�V�W�I�J�?�@�=�>�J�L�v�x�;O;�副I�J�C�C��犪   ��� ��� ��� ��� ���    zzz�111�444�FFF�FFF�VVV�ZZZ�PPP�ZZZ�ddd�^^^�___�ggg�nyn�n�o�\�]�N�O�V�W��à�      ����䋱s�t��މ?   ��� ��� ��� ��� ���    ����666�888�KKK�JJJ�ZZZ�___�UUU�___�lll�eee�fff�mmm�}}}�����r�s�d�e�������      ��� �����      ��� ��� ��� ��� ���    ����<<<�===�QQQ�MMM�^^^�ccc�XXX�eee�ttt�jjj�lll�rrr�����������������vvv�����      ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ����<<<�@@@�XXX�OOO�aaa�eee�\\\�jjj�{{{�qqq�rrr�www�����������������www�����      ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ����===�EEE�^^^�PPP�ccc�ggg�^^^�nnn�����www�xxx�~~~�������������������������      ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ����>>>�KKK�ddd�RRR�fff�jjj�___�sss�����|||�|||�����������������������������      ��� ��� ��� ��� ���             ���    ���dfff�bbb�{{{�eee�xxx�{{{�ppp�������������}}}����������������������������y      ��� ��� ��� ��� ���    �vh            ������r���У���������������������č��ʈ�����������ŷ������������������s���"   ��� ��� ��� ��� ��� ��� ��}���͞~eD         ��t(�Ju�t?���������~~~�KICp               cccq��������xxx�R      ��� ��� ��� ��� ��� ��� ��� ��~��s��[͑u^K   ��j8�N�� ��u;���������~~~�`U<z6)	      ���    cccq��������xxx�Q      ��� ��� ��� ��� ��� ��� ��� ��m��k ��m ��Zͽ�yq�O��z ��{ ��v7���������~~~�r^7��k0|sa
   ���    cccq��������xxx�Q      ��� ��� ��� ��� ��� ��� ��� �h��f ��j ��m ���/��s ��w ��x ��w5���������~~~��k=���\:            aaat��������xxx�   O      ��� ��� ��� ��� ��� ��� ��� �c��c ��f ��j ��m ��q ��s ��y��w,Ƭ�����������~te�   -            ^^^���������vvv�A      ��� ��� ��� ��� ��� ��� ��� �^��` ��c ��f ��j ��m ��u��x	��}�����������vvv�[[[�RRR�SSS�SSS�WWW�eee���������lll�   ,      ��� ��� ��� ��� ��� ��� ��� �Z��\ ��` ��c ��f ��o	��t��v	��Ѝ�}���������������������������������������������ddd�         ��� ��� ��� ��� ��� ��� ��� �U��Y ��\ ��` ��j��o��q��r	���"�հ������������������������������������������ggg�+++0      ��� ��� ��� ��� ��� ��� ��� ��� �Q��U ��Y ��e��l��m��n��p	��t��nԤ��{���蒒��������������xxx�uuu�mmm�eee�+++$   	   ��� ��� ��� ��� ��� ��� ��� ��� ��� �Xw�Z��`��h��i��j��k��l
��n��t	���jӴ��VZZZ            	      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ́[
�O��g��e��f��g��i��i
��j��m��o ���m�׭�5                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �f�Z��O��P��Q��S��U��V���W���a����o��|
   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���������������������  �  �  �  �  �  !�  s�  {�  �  �  �  �  �� �������� �� ��  �  �  �  ����������(   *   T                              ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                       ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                   "   $   &   (   *   ,   .   /   ,   $         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       �ܑ:�ꇶ}��|��{��{��z��z��z��y��y��{��s�|�5T8R   ,      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���xg�j��� � � � � � � � � � � � � � � � � � � � ������HtN\   "   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                     ����茯#�$� � � � � � � � � � � � � � � � � � � � ���J�K����   )   ��� ��� ��� ��� ��� ��� ��� ��� ���                                                 V�V�拰!�#� � � � � � � � � � � � � � � � ���=�=�C�C�����-   ��� ��� ��� ��� ��� ��� ���                                                          &:&�ሴ �"� � � � � � � � � � � � ���7�7�=�=�C�C�����*1   ��� ��� ��� ��� ��� ��� ���       	      #   ,   /   0   0   0   0   0   0   0   0   0   0   0   0   0   1:���	�	� � � � � � � � ���1�1�7�7�=�=�B�B����+0   ��� ��� ��� ��� ��� ���       DDD���Fuuu^jjjjhhhnhhhnjjjolllolllommmpmmmpoooqppprppprrrrrssssssssuuutwwwv�Ê�.�0� � � � � � � � ���,�,�2�2�7�7�=�=�B�B����-.   ��� ��� ��� ��� ��� ���       ���Mttt�]]]�ccc�mmm�mmm�hhh�^^^�ppp��������������������������������������;�<��� � � � � � ���&�&�,�,�1�1�7�7�<�<�B�B����/,   ��� ��� ��� ��� ��� ���       ����GGG��***�111�444�===�>>>�<<<�888�888�???�@@@�>>>�AAA�DDD�IJI�e{e�8�9������� � �
�
� � �&�&�,�,�1�1�6�6�<�<�B�B����1*   ��� ��� ��� ��� ��� ���       ����HHH��)))�000�333�===�AAA�@@@�<<<�===�EEE�FFF�DDD�FFF�JJJ�Zh[�=�>�&�'����������� � �&�&�+�+�1�1�6�6�<�<�A�A���� 3 (   ��� ��� ��� ��� ��� ���       ����LLL��+++�444�777�AAA�HHH�EEE�AAA�AAA�KKK�LLL�JJJ�KKK�PWP�BoC�6v7�2�3�+�,�� ���� � �!� � �%�%�+�+�0�0�6�6�<�<�A�A����"6"&   ��� ��� ��� ��� ��� ���       ����SSS�   �000�888�999�EEE�NNN�KKK�EEE�FFF�RRR�SSS�OOO�OQO�I^I�EiF�CuD�@�A�8�9�-�.�-�.�(�)�.�/�"�#�'�'�{�~�K�L�6�6�;�;�A�A����$:$#   ��� ��� ��� ��� ��� ���       ����NNN�"""�444�===�===�JJJ�RRR�PPP�III�JJJ�WWW�YYY�UUU�TTT�T\T�RhR�QuR�O�P�G�H�?�@�9�:�1�2�<�=�-�.�u�wۄƈB�银O�P�;�;�@�@����-H-   	��� ��� ��� ��� ��� ���       ����FFF�$$$�888�BBB�@@@�NNN�VVV�VVV�MMM�NNN�]]]�___�ZZZ�ZZZ�]]]�_g_�^t^�_�`�Y�Z�M�N�E�F�<�=�J�K�{�}�d�hE   V�V	�엶T�U�@�@���� 0    ��� ��� ��� ��� ��� ���       ����???�&&&�<<<�GGG�CCC�QQQ�ZZZ�ZZZ�PPP�QQQ�ccc�fff�___�___�bbb�hhh�nvn�q�q�j�k�Z�[�Q�R�G�H���������       	   ����혷a�c���      ��� ��� ��� ��� ��� ���       ����HHH�'''�@@@�KKK�DDD�TTT�]]]�___�TTT�UUU�iii�kkk�ccc�eee�eee�mmm�yyy�����~�~�i�j�`�a�o�p��������r      	   ��� �ے�񞽙�9   ��� ��� ��� ��� ��� ��� ���       ����QQQ�)))�EEE�PPP�FFF�WWW�aaa�aaa�WWW�WWW�nnn�qqq�iii�iii�jjj�qqq����������y�y�z�z�xzx��������q      	   ��� ��� ������ ��� ��� ��� ��� ��� ��� ��� ���       ����UUU�+++�HHH�TTT�GGG�YYY�ddd�ddd�YYY�ZZZ�ttt�www�nnn�nnn�ooo�vvv���������������������xxx��������q      	   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ����UUU�---�MMM�YYY�III�[[[�fff�eee�\\\�\\\�yyy�|||�rrr�sss�uuu�yyy���������������������zzz��������p      	   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ����WWW�...�PPP�```�KKK�^^^�iii�ggg�^^^�___�~~~�����vvv�vvv�xxx�}}}���������������������}}}��������n         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ����WWW�000�UUU�eee�LLL�___�jjj�ggg�^^^�aaa���������zzz�{{{�}}}�����������������������������󙙙i         ��� ��� ��� ��� ��� ��� ���          ��� ��� ���    ���zYYY�222�YYY�jjj�KKK�```�kkk�iii�]]]�bbb���������������������������������������|||�����\         ��� ��� ��� ��� ��� ���                   ���    ���>zzz�ZZZ�zzz�����jjj�}}}���������yyy�����������������rrr������������������������������������Ϳ��C   	   ��� ��� ��� ��� ��� ��� ���    +% 
                  ������D��������������������������������ǔ��Ώ��̏���������������ܺ��������������������������K���      ��� ��� ��� ��� ��� ��� ���    ����Ϥ�^         	         
ֲ�P֒)ovn_Բ�����������fee�   7      
               	eee�������������hhh�   C   "      ��� ��� ��� ��� ��� ��� ��� ��� ��� �{j��n���Yռ�ui            ߶�c�.��} uyn]ش�����������ffe�0! @      	      ���       eee�������������hhh�   B       	   ��� ��� ��� ��� ��� ��� ��� ��� ��� �g��)��o ���Yظ�sm   "   ޲�z�0��~ ��{ �|o\۵�����������ffe�W; LQ8 &('$   ��� ���       eee�������������hhh�   B       	   ��� ��� ��� ��� ��� ��� ��� ��� ��� �z�y��l ��n ��Yٵ�qoګ���1��z ��{ ��z �~oZ߷�����������ffe�tL X�Y3��h   ��� ���       eee�������������hhh�   A       	   ��� ��� ��� ��� ��� ��� ��� ��� ��� 變z�u��i ��k ��n ���Y��2��u ��w ��y ��y ��oY㹹����������ffe��Zd��TMnfY               eee�������������hhh�   A      	   ��� ��� ��� ��� ��� ��� ��� ��� ��� �{z�r��f ��i ��k ��n ��p ��s ��u ��w ��y��pX溺����������hgf���N�KC:1         	   	      ccc�������������hhh�   =         ��� ��� ��� ��� ��� ��� ��� ��� ��� �wz�p��c ��f ��i ��k ��n ��p ��s ��x��z��tQⰰ����������www�WSNw9   )   #   !   !   #   (bbbӗ�����������fff�   7         ��� ��� ��� ��� ��� ��� ��� ��� ��� �r{�m��a ��c ��f ��i ��k ��n ��t��y
��x�̀1͓���������������qqq�YYY�EEE�GGG�GGG�GGG�GGG�^^^�fff�������������ddd�   -      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �n{�j��^ ��a ��c ��f ��i ��p	��u��v
��z��ˀ~}���������������������www�vvv�vvv�vvv�vvv���������������������bbb�         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �j{�g��\ ��^ ��a ��c ��l
��r��r��t
��x��ֻ��諫������������������������������������������������������ccc�)         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �f{�d��Y ��\ ��^ ��i��n��o��p��q
��t���J�ܹ�����Ӧ�����������������������������������������������bbb�SSSe         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �bz�b��V ��Y ��e��k��l��m��n��o
��p��x���k�ή������|||񁁁�������������|||�rrr�ppp�jjj�eee�eee�!         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �e]�d��T ��`��h��j��j��k��k��l��n��p	��w���f�Ѭ��ddd1mmm&eee2kkk@iiiAeee?XXX=UUU<                  ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ތc�~C��]��f��f��g��h��h��i��j��k��l��n��r���]�߱�q                              ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �_}ۃK��e��d��e��f��g��g��h��h	��j��k��m���!���ز�(                  ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �bB�a��^��`��b��d��f��i���k���m���o���u����w�      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ������  ������  �����  �����  ���� �  ���� �  ���� �  ���� �  ���� �  ��   �  �    �  �    �  �    �  �    �  �    �  �   p�  �   x�  �   ��  �   ��  �   ��  �   ��  �   ��  �   ��  ��  ��  ��  ��  �� ��  �����  �����  � ���  � ���  � ���  � ��  � ���  �  ��  �  ��  �  ��  �  ��  �  ?��  �����  �����  � ����  �����  (   0   `                              ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���          
                   !   #   %   &   (   )   *   (   #            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ~˃9�ڈp|ׁ�x�~�v�|�u�z�s�{�s�z�q�x�p�w�o�v�n�u�n�u�[�aq&C   0         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���퓮e�i�;�=�1�3�1�3�1�4�1�4�1�4�1�4�1�4�1�4�1�4�1�4�3�6�Q�W����W�]s   /      	��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���씯*�,� � � � � � � � � � � � � � � � � � � � � � � � � � �������9_@P   !   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                 ���
�따*�,� � � � � � � � � � � � � � � � � � � � � � ���@�@�d�e�~ۅ�   %   ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                          VyV�鑳*�,� � � � � � � � � � � � � � � � � � ���;�;�A�A�K�K����   &   ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                +=+�⎹+�,� � � � � � � � � � � � � � ���6�6�<�<�@�@�E�E�����   %   ��� ��� ��� ��� ��� ��� ��� ���                '   ,   .   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   0 9����� � � � � � � � � � ���1�1�6�6�;�;�@�@�E�E�����   $   ��� ��� ��� ��� ��� ��� ��� ���       @@@$YYYDLLLTGGGZEEE]GGG]GGG]GGG]III^III^III^KKK_KKK_KKK_MMM_MMM_MMM_PPP`PPP`PPP`OOOa���S�U� � � � � � � � � � ���,�,�1�1�6�6�;�;�@�@�E�E�����   #   ��� ��� ��� ��� ��� ��� ���       ���+����|||�}}}��������􊊊�����yyy��������򦦦𦦦響��﨨�響��שּׁ����Ǳ�]�_��� � � � � � � � ���'�'�,�,�1�1�6�6�;�;�@�@�D�D�����   !   ��� ��� ��� ��� ��� ��� ���       ���Lhhh�...�***�333�777�;;;�AAA�BBB�BBB�>>>�???�@@@�CCC�CCC�BBB�EEE�GGG�KKK�OOO�gwh�N�P���	�
��� � � � �
�
�"�"�'�'�,�,�1�1�6�6�:�:�?�?�D�D�����      ��� ��� ��� ��� ��� ��� ���       ���Paaa��###�---�111�444�<<<�>>>�>>>�:::�999�<<<�BBB�CCC�AAA�CCC�EEE�JJJ�]h]�K�M�� �����	�
�������"�"�'�'�,�,�1�1�5�5�:�:�?�?�D�D�����      ��� ��� ��� ��� ��� ��� ���       ���Ohhh��###�---�111�444�>>>�CCC�DDD�>>>�>>>�@@@�HHH�HHH�FFF�GGG�KKK�W\W�I~J�-{.�)�*�"�#�����������"�"�'�'�,�,�0�0�5�5�:�:�?�?�D�D����      ��� ��� ��� ��� ��� ��� ���       ���Nooo��$$$�111�555�888�BBB�HHH�JJJ�BBB�AAA�EEE�MMM�NNN�KKK�KKK�MPM�GiH�:p;�8z9�3�4�,�-�"�#���#�$�#�$� �!�!�!�&�&�,�,�0�0�5�5�:�:�?�?�D�D�����      ��� ��� ��� ��� ��� ��� ���       ���Nuuu��'''�555�888�;;;�EEE�LLL�OOO�EEE�FFF�III�SSS�TTT�PPP�PPP�LZL�HeI�EnF�CyD�?�@�8�9�/�0�/�0�*�+�,�-�*�+�"�#�/�/����S�S�5�5�:�:�>�>�C�C����      ��� ��� ��� ��� ��� ��� ���       ���Mooo��)))�999�<<<�>>>�III�QQQ�TTT�JJJ�III�MMM�XXX�YYY�TTT�TTT�UYU�RcR�PmQ�PyQ�M�N�F�G�?�@�9�:�2�3�6�7�6�7�/�0��هلĈ<�혺V�W�9�9�>�>�C�C����      	��� ��� ��� ��� ��� ��� ���       ���Lddd��,,,�===�???�AAA�LLL�TTT�YYY�LLL�LLL�QQQ�]]]�^^^�YYY�YYY�ZZZ�^b^�\m\�]z^�[�\�V�W�J�K�D�E�;�<�A�B�H�I�΄�h�l;   ^�u�Z�[�>�>�D�E�����      ��� ��� ��� ��� ��� ��� ���       ���LXXX��...�BBB�CCC�CCC�OOO�XXX�___�PPP�PPP�UUU�ccc�ccc�]]]�^^^�^^^�eee�hlh�j{j�k�l�d�e�V�W�P�Q�D�E�O�P��̗�|�~a      	   �ȏ	��^�_�W�X���      ��� ��� ��� ��� ��� ��� ���       ���K[[[��111�FFF�FFF�DDD�RRR�ZZZ�bbb�SSS�RRR�WWW�iii�hhh�aaa�bbb�bbb�iii�ooo�z~z�{�{�t�u�c�d�\�]�P�Q���������cccN      	      ���򞽘����B      ��� ��� ��� ��� ��� ��� ���       ���Jhhh��333�JJJ�JJJ�FFF�UUU�]]]�eee�VVV�UUU�[[[�mmm�nnn�eee�fff�fff�mmm�ttt�������������q�r�j�k�s�s���������cccN      	   ��� ��� �����Z      ��� ��� ��� ��� ��� ��� ��� ���       ���Isss�!!!�555�NNN�MMM�HHH�WWW�___�ggg�XXX�WWW�^^^�rrr�sss�jjj�kkk�kkk�qqq�www�������������������yyy�yyy�����```M      	   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ���Ivvv�!!!�888�SSS�PPP�JJJ�YYY�aaa�jjj�[[[�YYY�aaa�www�xxx�nnn�nnn�nnn�uuu�{{{���������������������xxx�qqq�����```M      	   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ���Hvvv�"""�:::�XXX�TTT�KKK�[[[�ddd�lll�[[[�\\\�ccc�{{{�|||�rrr�rrr�rrr�yyy�~~~���������������������{{{�xxx�����aaaL      	   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ���Gvvv�"""�===�\\\�WWW�LLL�]]]�eee�nnn�ZZZ�^^^�fff������vvv�vvv�vvv�}}}�������������������������}}}���������bbbK         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ���Exxx�$$$�@@@�```�[[[�MMM�]]]�hhh�ppp�[[[�___�hhh���������yyy�zzz�zzz��������������������������������������fffF         ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��� ��� ���       ���Axxx�&&&�CCC�eee�___�MMM�```�jjj�sss�ZZZ�aaa�jjj���������}}}�~~~�~~~�����������������������������}}}���������uuu=         ��� ��� ��� ��� ��� ��� ���                   ��� ���    ���:����+++�FFF�jjj�bbb�MMM�aaa�jjj�sss�ZZZ�```�lll�������������������������������������������������{{{�������Ʀ���0   
   ��� ��� ��� ��� ��� ��� ��� ���             	         ���    ���#������������������������������������������������񴴴򓓓�zzz�yyy����������������������������������������gEEE      ��� ��� ��� ��� ��� ��� ��� ���    �|lp`T         	         %%%����¯Uհu~~}|�����������������xxx����J���:���3���0���1���2���2���4���<�����������������sssx���U���>���      ��� ��� ��� ��� ��� ��� ��� ��� ���    ��������LA9)         
         ϰ�D�L|�x gjif�������������nnn�MLG�   %                        eee�������������ggg�Y   *         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �����q��~���@700            Բ�S�Q�� z�x ujif�������������nnn�YSD� )            ���          eee�������������ggg�X   )         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� 湝F��A��n ��~��?5.2       ҭ�d�T��~ ��~ ��x �kif�������������nnn�eY@�S9 4C1      ��� ��� ���       fff�������������ggg�X   )         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� 깛N��6��l ��m ��~��<3,5ˣ�x�W��z ��{ ��| ��y �kif�������������nnn�n^>�wP @�e#��w   ��� ��� ���       ggg�������������ggg�X   )         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� 贕O��5��i ��l ��m ��~����Z��v ��x ��y ��z ��x �lie�������������nnn�xb;��bM��h9_[T	                  hhh�������������ggg�W   (         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� 豑O��3��f ��i ��k ��m ��u��r ��s ��u ��x ��x ��y�lie�������������nnn��g;���^iMH@   
               	   ggg�������������ggg�V   &         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� 欌P�2��d ��f ��i ��k ��m ��o ��r ��s ��u ��z��y�lid�������������uuu���f�3/)A   #                     !ccc�������������ggg�N   #      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� 橇P�~0��b ��d ��f ��i ��k ��m ��o ��r ��w��z	��y�}sh�����������������oon�M   :   1   -   ,   ,   -   0111Xjjj�������������ccc�   :         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� 䤂Q�z/��` ��b ��d ��f ��i ��k ��m ��t��x��x	��}ƚ~b꯯��������������www�nnn�\\\�[[[�[[[�[[[�[[[�[[[�aaa�bbb�����������������bbb�   0         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �~Q�x-��] ��` ��b ��d ��f ��i ��q
��t��u��w	���ц=ւ���������������������������|||�|||�|||�|||�{{{���������������������{{{�aaa�   #         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �yQ�v,��[ ��] ��` ��b ��d ��l��r��s��s��u
��~��+՜�������������������������������������������������������������������bbb�,         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �uQ�r*��Y ��[ ��] ��` ��j��o��o��q��q��r	��z����毟�r������������������������������������������������������������bbb�UUUo      
      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �rP�p)��V ��Y ��[ ��f��m��m��m��n��o��p	��v���0��֏��Y���ˀ���������������������������������������xxx�fff�bbb�CCC9      
      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �pK�o*��T ��V ��c��j��j��k��l��l��m��n	��q	��w���/��և�{MzzzG�uuu�lll�kkk�jjj�hhh�eee�ccc�eee�eee�LLL<               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ݍe!�~B��R ��`��g��h��h��i��j��k��k��l	��m��q��v���'�����}rl9RRR+++      
   
   
   
   
   
   	               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �`��b��e��e��f��g��g��h��i��i��j
��j��l��n��o�������ʁk\                                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �h#�g��x;��g��d��d��f��f��f��h��h
��i��i��k��m��}����� e      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �}X	�en�g��i��l��o���q���t���w���y���|����������������綗.      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ������  ������  ���� ?  ����   ����   ����   ����   ����   ����   ����   ��     ��     ��     ��     ��     ��     ��    ��  �  ��  �  ��  �  ��  �  ��  �  ��  �  ��  �  ��  �  ��  �  ��  �  ��  �  ��  �  ����  ����  ����  ����  � ��  � ��  � ��  � ��  � ��  �   �  �   �  �   ��  � ��  � ��  � ���  � ���  � ?���  � ?���  � ���  (   @   �                              ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                       
                                                   	             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                               !   !                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                             "   $   &   (   )   +   ,   .   /   1   2   3   3   3   /   *   !            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���           QqQ�ێS�蓇�葤�䎧�ጩ�ߋ������ߊ��݋��܊��ۉ��ډ��و��؈��ه�؆�~ԇ�n�u�AjF^   ;   1   #         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���        ��<����y�~�U�Y�E�H�E�H�E�H�E�H�E�H�E�H�E�H�E�I�E�I�E�I�E�I�E�I�E�I�E�I�H�M�h�o�����ڇ�+G   0         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���     �ի����e�h� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���n�t����:   '      
��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                �߫��N�Q� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���B�B�����s�z�   ,      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                              �ѡ��O�Q� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���>�>�C�C�h�k����   /      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                   �����O�Q� � � � � � � � � � � � � � � � � � � � � � � � � � ���:�:�?�?�B�B�P�P�����   /      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                    
                                                                     ZvZ�O�R� � � � � � � � � � � � � � � � � � � � � � ���6�6�;�;�?�?�B�B�F�F�����   /      ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                               :K:,���O�R� � � � � � � � � � � � � � � � � � ���2�2�7�7�;�;�>�>�B�B�F�F�����   .      ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                        )   .   1   2   2   2   2   2   2   2   2   2   2   2   2   2   2   2   2   2   2   2   2   3   3   57O7J���-�/� � � � � � � � � � � � � � ���/�/�3�3�7�7�;�;�>�>�B�B�F�F�����   ,      ��� ��� ��� ��� ��� ��� ��� ��� ��� ���          	   #3>F


I


J


J


J


J


J


J


J


J


J


J


J


J


J


J


J


J


J


J


J


J


J


K"R�̋�R�U��� � � � � � � � � � � � ���+�+�0�0�3�3�7�7�:�:�>�>�B�B�E�E�����   +      ��� ��� ��� ��� ��� ��� ��� ��� ���           """���F���o���������������������������������������������������������������������������������������������������������٬�S�V��� � � � � � � � � � � � ���'�'�,�,�/�/�3�3�7�7�:�:�>�>�B�B�E�E�����   *      ��� ��� ��� ��� ��� ��� ��� ��� ���           ���-���innn�^^^�\\\�ccc�iii�nnn�lll�hhh�aaa�WWW�ggg�sss����������������������������������������������������������X�Z����� � � � � � � � � � �
�
�#�#�(�(�,�,�/�/�3�3�6�6�:�:�>�>�A�A�E�E�����   )      ��� ��� ��� ��� ��� ��� ��� ��� ���           ���D����MMM��###�***�111�222�555�;;;�>>>�???�???�:::�999�888�888�===�===�>>>�<<<�===�@@@�BBB�EEE�GGG�NNN�s�t�L�M�����	�
��� � � � � � �	�	���$�$�(�(�+�+�/�/�3�3�6�6�:�:�>�>�A�A�E�E�����   '      ��� ��� ��� ��� ��� ��� ��� ��� ���           ���Fyyy�CCC��"""�)))�111�111�333�:::�>>>�>>>�>>>�:::�999�999�:::�AAA�BBB�BBB�@@@�AAA�DDD�FFF�III�NNN�k~l�L�M���������	�
��� � ����� � �$�$�(�(�+�+�/�/�2�2�6�6�:�:�=�=�A�A�E�E�����   &      ��� ��� ��� ��� ��� ��� ��� ��� ���           ���F}}}�FFF��"""�)))�111�000�222�:::�???�AAA�BBB�>>>�<<<�===�===�EEE�FFF�FFF�CCC�DDD�GGG�III�MMM�ana�J�K�)}*�%�&�!�"�������	�
������� � �#�#�'�'�+�+�/�/�2�2�6�6�:�:�=�=�A�A�D�D�����   %      ��� ��� ��� ��� ��� ��� ��� ��� ���           ���E����HHH��"""�)))�222�222�444�===�BBB�EEE�GGG�AAA�???�???�@@@�III�JJJ�KKK�HHH�HHH�JJJ�MMM�XaX�GxH�2t3�1|2�-�.�)�*�"�#������������� � �#�#�'�'�+�+�.�.�2�2�6�6�9�9�=�=�A�A�D�D�����   #      ��� ��� ��� ��� ��� ��� ��� ��� ���           ���E����JJJ��$$$�,,,�666�444�777�@@@�EEE�III�KKK�DDD�BBB�BBB�CCC�MMM�NNN�OOO�KKK�KKK�MMM�MRM�GiH�<l=�:s;�9{:�6�7�1�2�*�+�"�#� �!�$�%�#�$�$�%�"�#���#�#�'�'�,�,�.�.�2�2�6�6�9�9�=�=�@�@�D�D�����   !      
��� ��� ��� ��� ��� ��� ��� ��� ���           ���D����NNN��&&&�///�999�777�999�CCC�HHH�MMM�OOO�GGG�EEE�EEE�FFF�QQQ�SSS�SSS�OOO�OOO�PRP�J\J�FcG�DjE�CsD�AzB�?�@�:�;�2�3�-�.�0�1�+�,�(�)�,�-�+�,�#�$�#�#�)�)�߃�o�r�2�2�5�5�9�9�=�=�@�@�D�D�����         	��� ��� ��� ��� ��� ��� ��� ��� ���           ���D����MMM��'''�222�===�:::�<<<�EEE�KKK�PPP�SSS�JJJ�HHH�HHH�III�UUU�WWW�WWW�RRR�RRR�RSR�P[P�PdP�LiM�KqL�JzK�H�I�D�E�<�=�:�;�7�8�1�2�-�.�4�5�3�4�(�)�'�'�y�{�ꠡ���q�t�5�5�9�9�<�<�@�@�D�D�����         ��� ��� ��� ��� ��� ��� ��� ��� ���           ���C����HHH��)))�444�@@@�<<<�===�HHH�MMM�SSS�WWW�MMM�JJJ�KKK�KKK�YYY�ZZZ�[[[�VVV�WWW�VVV�XYX�XcX�ThT�TqU�U{V�S�T�P�Q�H�I�A�B�?�@�8�9�4�5�<�=�<�=�0�0�s�u�ޜ�+v�v����t�v�8�8�<�<�@�@�D�D�����         ��� ��� ��� ��� ��� ��� ��� ��� ���           ���Czzz�DDD��+++�777�DDD�???�???�JJJ�PPP�UUU�[[[�QQQ�MMM�MMM�MMM�]]]�___�___�YYY�YYY�YYY�[[[�`a`�\g\�]q]�_|`�^�_�[�\�Q�R�K�L�G�H�?�@�;�<�E�F�G�H�w�y�ʔ�      �ɏ����v�x�<�<�@�@�F�G�����      
   ��� ��� ��� ��� ��� ��� ��� ��� ���           ���Bqqq�@@@��---�:::�GGG�AAA�@@@�LLL�RRR�XXX�^^^�SSS�OOO�OOO�PPP�aaa�bbb�ccc�]]]�^^^�]]]�^^^�ddd�fgf�grg�j~j�i�j�g�h�Z�[�T�U�P�Q�F�G�B�C�N�O��ȃ��ͫ�-      	      ������x�z�@�@�Z�[�����         ��� ��� ��� ��� ��� ��� ��� ��� ���           ���Bmmm�@@@��...�===�KKK�DDD�BBB�NNN�SSS�ZZZ�aaa�VVV�RRR�QQQ�SSS�eee�fff�ggg�```�```�```�aaa�ggg�iii�pqp�v�v�v�v�s�t�f�g�]�^�X�Y�N�O�J�K�z�|��κ圞�x   *      	         ������{�~��������         ��� ��� ��� ��� ��� ��� ��� ��� ���           ���Avvv�DDD��111�???�OOO�FFF�CCC�OOO�VVV�\\\�bbb�XXX�TTT�SSS�TTT�hhh�jjj�kkk�ccc�ccc�ddd�ddd�jjj�mmm�ttt�������������s�t�g�h�b�c�W�X�k�l��������ۜ��w   *      	             �����Ȥ���ێ         ��� ��� ��� ��� ��� ��� ��� ��� ���           ���A}}}�III�   �111�BBB�SSS�HHH�EEE�RRR�XXX�^^^�eee�[[[�UUU�UUU�VVV�kkk�nnn�nnn�fff�ggg�ggg�fff�mmm�ppp�xxx���������������r�s�m�n�m�n����������ޛ��w   *      	      ���         �����:              ��� ��� ��� ��� ��� ��� ��� ��� ���           ���@����OOO�!!!�444�EEE�VVV�III�EEE�TTT�ZZZ�```�hhh�]]]�WWW�XXX�XXX�ppp�qqq�rrr�iii�jjj�kkk�jjj�ppp�sss�{{{�����������������|�|�|�|���vvv�|||����ᛛ�w   *      	      ��� ��� ���                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���           ���@����PPP�!!!�555�HHH�ZZZ�LLL�FFF�TTT�[[[�bbb�jjj�^^^�YYY�YYY�[[[�rrr�uuu�vvv�mmm�mmm�mmm�lll�sss�uuu��������������������������|||�www�ttt����䚚�v   *      	      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���           ���@����QQQ�###�777�JJJ�___�NNN�GGG�VVV�]]]�ddd�jjj�^^^�[[[�ZZZ�\\\�vvv�yyy�yyy�ooo�ppp�ppp�ppp�vvv�xxx������������������������������xxx�nnn����皚�v   *      	      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���           ���@����QQQ�"""�999�MMM�ccc�PPP�HHH�YYY�___�fff�mmm�___�]]]�]]]�]]]�yyy�|||�}}}�rrr�sss�sss�sss�yyy�zzz���������������������������������{{{�xxx����晙�t   )      	      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���           ���@����RRR�###�;;;�PPP�ggg�RRR�HHH�YYY�```�ggg�ooo�___�]]]�]]]�___�|||���������vvv�vvv�vvv�uuu�|||�|||���������������������������������|||��������⚚�t   (            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���           ���=����SSS�$$$�===�RRR�kkk�TTT�III�[[[�aaa�iii�ppp�```�]]]�___�___�������������xxx�yyy�yyy�yyy�����������������������������������������~~~��������ݛ��q   &            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���           ���;����SSS�%%%�???�UUU�ppp�VVV�III�[[[�ccc�jjj�qqq�```�^^^�aaa�bbb�������������zzz�{{{�{{{�{{{�������������������������������������������������آ��l   "             ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                      ��� ���           ���8����TTT�'''�AAA�XXX�ttt�YYY�III�\\\�ccc�jjj�sss�```�\\\�aaa�ccc�������������}}}�~~~�������������������������������������������|||��������ѭ��d                ��� ��� ��� ��� ��� ��� ��� ��� ���                                        ���6����^^^�(((�DDD�[[[�yyy�ZZZ�III�]]]�eee�lll�sss�aaa�\\\�```�ccc������������������������������������������������������������������zzz�������ü���[      	      ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                      ���%���Y����aaa�nnn�������������qqq�������������������������������������������������yyy�nnn�zzz����������������������������������������������������z���?             ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                   
                  ������@���\�������ݠ��𞞞������������������������㵵�к����������������������ů��Π��ԑ��ܒ��ۢ��թ��𳳳������������������������ݼ����������y���^{{{             ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ɫ�7            	                  	���"�ūd׫f}��l�xxx�����������������rrr�mmm�___F~~~7���+���&���$���#���#���#���$���$���&���+~~~�������������������ppp�ccc~dddR���?���*   
             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��}�˦�����
            	            	&"���a�J~�z f�rU�kkk�����������������bbb�RPM�   /                                 ggg�ttt�����������������\\\�000j   6   !                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �Þ���4���_�给�	%               
   )%!�ßp�N�ـ s�z p�sS�kkk�����������������bbb�ZUK� 3                                   	hhh�vvv�����������������\\\�000j   6                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �Ǣ��o��p ���_�乗�
	(             �Þ��O�� ��~ ~�y z�tQ�kkk�����������������bbb�`YH�<* ;'                  ��� ���          	hhh�www�����������������\\\�000j   5                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �xe�����l ��n ��p ���_�㸗�
	)   "   �����P��~ ��~ ��} ��y ��tP�kkk�����������������bbb�h]F�W; DV< )D0             ��� ���          	hhh�yyy�����������������\\\�000j   5                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��s�����k ��l ��n ��o ���`�ⷖ�
,*罚��Q��z ��{ ��| ��| ��y ��tN�kkk�����������������bbb�n`E�oK LwQ 1�^	��x          ��� ���          	hhh�{{{�����������������\\\�000j   5                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��l�����h ��j ��k ��m ��o ���`�ⷖ�滙��S��w ��y ��y ��z ��z ��y ��uM�kkk�����������������bbb�tbC��U S�a:��Z4���                           	ggg�}}}�����������������\\\�000i   5                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��j�����f ��h ��j ��k ��m ��o ���`���T��t ��u ��w ��x ��x ��y ��x ��uL�kkk�����������������bbb�ydA��\ \��TW���-                        ggg�{{{�����������������\\\�111h   4                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �g�����e ��f ��h ��j ��k ��m ��o ��q ��s ��s ��u ��w ��x ��x ��z��vK�kkk�����������������bbb�~f?���P|��vJ                        
   fff�ttt�����������������\\\�111h   2                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �}e�����c ��e ��f ��h ��j ��k ��m ��o ��q ��r ��s ��u ��v ��{��z��uI�kkk�����������������eee��a}ik   ,                              eee�nnn�����������������\\\�222e   /                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �w_��~��a ��c ��e ��f ��h ��j ��k ��m ��o ��q ��r ��s ��y��{��z��w3�fff�����������������sss�yvr�K   :   .   '   #   "   !   !   "   #   &   -ccc�sss�����������������]]]�E   +      
      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �u]��{��` ��a ��c ��e ��f ��h ��j ��k ��m ��o ��q ��v��y
��z��{
���jii���������������������nnn�***`N   B   <   9   8   8   8   8   9   <K___���������������������aaa�   :   %             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �s[��x��^ ��` ��a ��c ��e ��f ��h ��j ��k ��m ��t	��x��x
��x	��}���usq���������������������www�lll�kkk�```�___�```�```�```�```�```�```�bbb�^^^�nnn�����������������zzz�bbb�   2                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �nV��u��\ ��^ ��` ��a ��c ��e ��f ��h ��j ��q
��u��v��w
��x��~��ʉ}q�����������������������������}}}�rrr�nnn�nnn�nnn�nnn�nnn�nnn�nnn�uuu�������������������������ccc�^^^�   (      
      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �lS��r��Z ��\ ��^ ��` ��a ��c ��e ��f ��n��s��s��t��u
��x��~�����6�~}|�������������������������������������������������������������������������������������xxx�aaa�   -               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �jQ��o��Y ��Z ��\ ��^ ��` ��a ��c ��l��p��q��r��r��s
��v��}�� ����Ღ�ؕ�����������������������������������������������������������������������������������^^^�HHHc         	          ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �iO��l��W ��Y ��Z ��\ ��^ ��` ��i��n��o��o��p��q��q
��t��z���N��ϳ�~~}T���ۘ�����������������������������������������������������������������������vvv�^^^�bbb�         
          ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �oS�i��U ��W ��Y ��Z ��\ ��g��m��m��m��n��n��o��p
��q
��w��}���w��Ī��T����������������������������������������������������������������yyy�ccc�bbb�MMMV         
             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �rT�g��S ��U ��W ��Y ��d��j��k��l��l��l��m��m��n
��o	��r��x��~���w��ũ�xwwL���M����{{{�rrr�ggg�^^^�\\\�\\\�\\\�\\\�\\\�\\\�\\\�^^^�bbb�eee�eee�                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� uL7��j��R ��S ��U ��b��i��i��i��j��k��k��l��l��l��m	��n��r��x��|���s��ŧ�mkj?jjj5lll-ddd$HHH""""""""""""                                        ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��jݿT��R ��`��g��g��h��h��h��i��j��j��k��l��k	��l��n��q
��v��y���m��ä�[ZX,RRR>>>      	                                                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �f~�{>��^��e��e��f��f��g��g��h��h��i��i��j��k	��k��k��n��o��q��u���h��ģ�0,*                                                    ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    f@-��l��~E��d��d��d��e��e��f��f��g��g��h��h��i
��j��j��k��m��m��o ��q ���y��Ȧ�                                                       ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���        у]��j��k���P��|=��|<��|;��}:��~:��9��8��8��8��7��7���6���6���5���5���K���z��Ü�ߵ�)             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���           �f#��pZ��m��o��q��t���v���y���{���~��������������������������������j칙5                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �����������������������������  �����  �����  �����  �����  �����  ������ ������ ������ ������ ��     ��     ��     ��     ��     ��     ��     ��     ��     ��    ��    ��    ?��    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ����   ��������������������������� ����� ����  ����  ����  ����  ����  ����  ����    ���    ���    ���    ?���   ?���   ����  ���� ������ ������  ������  �����  ������ �����(   �                                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                	   	   	   
   
   
   
                                                                        
   	                            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                    	                                                                                                               	                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                 
                                                                                                                           	                   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                                  !   !   "   "   #   #   $   $   %   %   %   %   $   #   "                         	               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                              
                               !   "   #   #   $   %   %   &   &   '   (   (   )   *   *   +   ,   ,   -   .   .   /   /   /   .   -   ,   *   '   #                  
            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                               	                         "   $   %   '   (   )   *   +   ,   ,   -   .   /   /   0   1   2   3   3   4   5   6   6   7   8   8   8   8   7   6   3   0   ,   (   "               	         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                              
         1S7%X�\:T�X=P�T?M{QBKxODIuMFHtLFGrKGFpIIEnHJDmHKDmHKClGLCkFMBiEMAhDN@gDO@fCP?eBQ>dAR>cAS>cAS<a?T<`?U<`?U;_>V;^=W:]=X:]=X0J   @   ?   >   <   9   5   0   *   $                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                           ~Ƅ+��x�������ܝ������������������������������������������������������������������������������������������������������������������������������ݒ�u�|�CnHd   A   =   8   1   +   #            
      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                      @`@���m��������������������������������������������������������������������������������������������������������������������������������������������������������}ʄ�H   ?   8   1   )   !            	   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���               ��+�����������^�b�3�5��� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���7�;�_�f������������JwOg   >   7   /   &            
   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���        �������������#�%� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �"�$�������������BjE`   ;   3   *   !            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���            ���<���Ǔ��M�O� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��������������A   7   .   $            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���           ���=���Ȕ��L�O� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �
�
�<�<�I�I���������yƃ�   :   0   '            	��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���               ���=���Ȕ��L�O� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �
�
�:�:�B�B�D�D�b�d���������6Y9Q   2   (            
��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                                                                                                                    ���=���ɔ��L�O� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �	�	�8�8�@�@�B�B�D�D�F�F���������l�t�   3   *             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                                                                                             ��@���ɔ��M�O� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �	�	�6�6�>�>�@�@�B�B�D�D�E�E�z�}������Ս�   4   *   !         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                                                                                                     ��A���˔��M�O� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �	�	�5�5�<�<�>�>�@�@�B�B�C�C�E�E�b�d��������   4   +   !         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                                                                                                              ��C���˔��M�O� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���3�3�:�:�<�<�>�>�@�@�B�B�C�C�E�E�L�L���������   4   +   !         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                      	   	   	   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
         �؛G���͔��M�O� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���1�1�8�8�:�:�<�<�>�>�@�@�A�A�C�C�E�E�G�G���������   4   *   !         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                             	                                                                                                                                                         �˒K���ϔ��M�P� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���0�0�6�6�8�8�:�:�<�<�>�>�@�@�A�A�C�C�E�E�G�G���������   3   *   !         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                           	                                                                                                                                                                  ���Q���є��M�P� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���.�.�4�4�6�6�8�8�:�:�<�<�>�>�?�?�A�A�C�C�E�E�G�G���������   3   *   !         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                       	                               !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   "   #   #   %v�|[���ӓ��M�P� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���,�,�2�2�4�4�6�6�8�8�:�:�<�<�>�>�?�?�A�A�C�C�E�E�G�G���������   2   )             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                        	                  #   &   (   *   +   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   -   -   .   /   1k�pd��ה��M�P� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���*�*�1�1�2�2�4�4�6�6�8�8�:�:�<�<�=�=�?�?�A�A�C�C�E�E�F�F���������   1   (             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                    	               #   (   -   0   3   5   6   7   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   9   9   :   ;FdIW��˔��b�e��� � � � � � � � � � � � � � � � � � � � � � � � � � � � ���)�)�/�/�1�1�2�2�4�4�6�6�8�8�:�:�<�<�=�=�?�?�A�A�C�C�E�E�F�F���������   1   (            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                $   +   1   7   ;   >   @   A   B   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   D   D   D   D   E?XB]�ߥÐ��]�`��� � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�'�-�-�/�/�0�0�2�2�4�4�6�6�8�8�:�:�;�;�=�=�?�?�A�A�C�C�D�D�F�F���������   0   '            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	         "&&&1###9!!!@FJNPRSSSSSSSSSSSSSSSSSSSTTTTTTTTTTTTTTTTTTTTTTTTUUUL]Li�ڥ����Y�[��� � � � � � � � � � � � � � � � � � � � � � � � � � � � ���%�%�+�+�-�-�/�/�0�0�2�2�4�4�6�6�8�8�:�:�;�;�=�=�?�?�A�A�C�C�D�D�F�F���������   /   '            
��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                    
   WWW ���Q���k���v���|������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������אߔ�V�X��� � � � � � � � � � � � � � � � � � � � � � � � � � � � ���#�#�)�)�+�+�-�-�.�.�0�0�2�2�4�4�6�6�8�8�9�9�;�;�=�=�?�?�A�A�B�B�D�D�F�F���������   .   &            
��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                    ��� ���a���k���r���|�������ڊ��݌��ގ��ݒ��ޔ��ݗ��ܙ��ܖ��ۖ��ܕ��ݔ��ޓ��ߑ������⍍�㑑�����ߘ��ݛ��ܞ��ڡ��ئ��֧��ԧ��է��է��ԩ��ԩ��Ԫ��ө��ө��ԩ��ԩ��ԩ��ԩ��ԩ��Ԫ��ԫ��ԫ��ԫ��Ԭ��ԭ��ԭ��Ԯ��ӯ��ӯ��ӱ��Բ��Գ��Է��ڿ���ܕ�X�Z�	�
��� � � � � � � � � � � � � � � � � � � � � � � � � � ���!�!�'�'�)�)�+�+�-�-�.�.�0�0�2�2�4�4�6�6�8�8�9�9�;�;�=�=�?�?�A�A�B�B�D�D�F�F���������   -   %            
��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 ���S���f���m����hhh�ccc�fff�jjj�mmm�qqq�uuu�yyy�|||������}}}�zzz�www�sss�lll�fff�^^^�ccc�mmm�vvv���������������������������������������������������������������������������������������������������������������������������׿��֓�Z�\��������� � � � � � � � � � � � � � � � � � � � � � ��� � �%�%�'�'�)�)�+�+�,�,�.�.�0�0�2�2�4�4�6�6�7�7�9�9�;�;�=�=�?�?�@�@�B�B�D�D�F�F���������   -   %            
��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 ������a���f����\\\�[[[�]]]�LLL�KKK�NNN�PPP�TTT�WWW�YYY�\\\�\\\�\\\�[[[�\\\�[[[�ZZZ�YYY�UUU�UUU�YYY�___�bbb�ccc�fff�iii�lll�nnn�nnn�nnn�rrr�rrr�rrr�rrr�rrr�qqq�ppp�qqq�qqq�rrr�sss�ttt�uuu�uuu�www�xxx�yyy�zzz�|||�}}}�~~~����������Ƈ�V�W�������	�
����� � � � � � � � � � � � � � � � � � �����#�#�%�%�'�'�)�)�+�+�,�,�.�.�0�0�2�2�4�4�6�6�7�7�9�9�;�;�=�=�>�>�@�@�B�B�D�D�F�F���������   ,   $            
��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���+���a���gmmm�UUU�JJJ���!!!�%%%�'''�,,,�000�222�333�000�333�666�:::�===�???�>>>�???�>>>�???�???�<<<�999�999�999�888�888�888�888�<<<�===�===�===�===�<<<�:::�;;;�<<<�===�???�@@@�@@@�AAA�DDD�EEE�EEE�GGG�JJJ�KKK�WZW�����u�v�P�R����������	������� � � � � � � � � � � � � � �����!�!�#�#�%�%�'�'�)�)�*�*�,�,�.�.�0�0�2�2�4�4�5�5�7�7�9�9�;�;�=�=�>�>�@�@�B�B�D�D�F�F���������   +   #            	��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���.���a���gddd�[[[�(((���!!!�%%%�'''�,,,�///�111�333�000�222�666�:::�<<<�>>>�>>>�>>>�>>>�???�???�<<<�999�999�888�888�777�777�777�===�>>>�>>>�???�???�???�===�===�>>>�???�@@@�AAA�CCC�CCC�EEE�GGG�HHH�III�LLL�VXV����q�s�N�P�������������	�
������� � � � � � � � � � �������!�!�#�#�%�%�'�'�)�)�*�*�,�,�.�.�0�0�2�2�4�4�5�5�7�7�9�9�;�;�<�<�>�>�@�@�B�B�D�D�F�F���������   *   #            	��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���-���a���gddd�___����   �$$$�'''�,,,�///�111�222�///�222�555�999�;;;�===�>>>�>>>�???�>>>�>>>�;;;�888�888�999�888�888�999�999�???�@@@�AAA�AAA�AAA�AAA�???�???�@@@�AAA�BBB�CCC�EEE�EEE�HHH�HHH�JJJ�LLL�VWV�z�z�m�n�N�O�����������������	�
������� � � � � � ���������!�!�#�#�%�%�'�'�(�(�*�*�,�,�.�.�0�0�2�2�3�3�5�5�7�7�9�9�;�;�<�<�>�>�@�@�B�B�D�D�F�F���������   *   #            	��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���.���`���ghhh�bbb����   �$$$�&&&�,,,�///�111�222�///�111�555�999�;;;�===�>>>�>>>�>>>�>>>�???�<<<�999�999�:::�:::�:::�:::�;;;�AAA�BBB�CCC�DDD�CCC�CCC�@@@�AAA�AAA�CCC�DDD�EEE�FFF�GGG�III�KKK�LLL�TUT�t}u�g�h�L�M�$�%� �!�� ���������������	�
������� � �����������!�!�#�#�%�%�'�'�(�(�*�*�,�,�.�.�0�0�2�2�3�3�5�5�7�7�9�9�:�:�<�<�>�>�@�@�B�B�D�D�F�F���������   )   "            	��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���.���`���glll�fff����   �$$$�&&&�,,,�///�111�222�...�111�444�888�:::�===�???�???�@@@�AAA�AAA�>>>�;;;�;;;�;;;�;;;�<<<�<<<�<<<�CCC�DDD�EEE�EEE�EEE�EEE�BBB�BBB�CCC�DDD�EEE�GGG�HHH�III�KKK�MMM�RSR�nsn�b�c�J�K�(|)�&~'�$�%�#�$�!�"���������������	�
�����������������!�!�#�#�%�%�&�&�(�(�*�*�,�,�.�.�0�0�1�1�3�3�5�5�7�7�9�9�:�:�<�<�>�>�@�@�B�B�D�D�E�E���������   (   !            	��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���.���`���gppp�hhh����   �$$$�&&&�,,,�///�111�222�...�000�555�888�<<<�>>>�AAA�BBB�BBB�CCC�DDD�@@@�===�>>>�===�===�===�>>>�>>>�EEE�FFF�GGG�GGG�GGG�GGG�EEE�EEE�EEE�EEE�GGG�HHH�III�KKK�MMM�RSR�hkh�\�]�I�J�-x.�+{,�*~+�'(�'�(�$�%�"�#���������������	�
�	�
�������������!�!�#�#�%�%�&�&�(�(�*�*�,�,�.�.�0�0�1�1�3�3�5�5�7�7�8�8�:�:�<�<�>�>�@�@�B�B�D�D�E�E���������   (   !            	��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���.���`���fuuu�mmm�����###�&&&�---�000�222�333�///�222�555�:::�===�???�BBB�DDD�EEE�FFF�FFF�BBB�>>>�???�???�???�>>>�???�???�GGG�HHH�III�III�JJJ�III�GGG�GGG�GGG�GGG�III�III�KKK�LLL�RRR�bdb�WzX�H�I�3t4�0w1�/z0�/0�+,�+�,�(�)�&�'�"�#�����������������������������!�!�#�#�$�$�&�&�(�(�*�*�,�,�.�.�/�/�1�1�3�3�5�5�7�7�8�8�:�:�<�<�>�>�@�@�B�B�C�C�E�E���������   '                	��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���.���_���fxxx�ppp����   �$$$�&&&�...�222�444�555�000�333�888�<<<�???�AAA�DDD�EEE�GGG�GGG�GGG�DDD�@@@�@@@�@@@�@@@�@@@�AAA�AAA�III�KKK�KKK�KKK�LLL�KKK�III�HHH�JJJ�III�JJJ�LLL�MMM�NNN�Z[Z�RqS�FxG�6o7�5s6�3u4�3z4�2}3�/0�/�0�,�-�*�+�&�'�!�"�������������������� �������!�!�"�"�$�$�&�&�(�(�*�*�,�,�.�.�/�/�1�1�3�3�5�5�6�6�8�8�:�:�<�<�>�>�@�@�B�B�C�C�E�E���������   &               	��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���.���_���f}}}�ttt����   �%%%�(((�///�333�666�777�111�444�888�===�@@@�CCC�EEE�HHH�HHH�III�JJJ�EEE�AAA�BBB�BBB�AAA�BBB�BBB�CCC�LLL�MMM�MMM�NNN�MMM�NNN�JJJ�JJJ�JJJ�JJJ�KKK�MMM�NNN�STS�LeM�DnE�;k<�9n:�9r:�7u8�7y8�7~8�3~4�3�4�1�2�.�/�*�+�%�&�"�#�� �����#�$�"�#�!�"� �!�� �#�$�"�#�����!�!�"�"�$�$�&�&�(�(�*�*�,�,�-�-�/�/�1�1�3�3�5�5�6�6�8�8�:�:�<�<�>�>�@�@�A�A�C�C�E�E���������   %               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���-���_���e����xxx����!!!�&&&�)))�111�555�777�888�222�666�:::�???�AAA�DDD�GGG�JJJ�KKK�KKK�KKK�GGG�CCC�CCC�CCC�CCC�DDD�DDD�EEE�MMM�OOO�OOO�OOO�OOO�OOO�LLL�MMM�LLL�LLL�MMM�NNN�PPP�G[G�DfE�@fA�>i?�=m>�=r>�;t<�;y<�;}<�89�8�9�5�6�2�3�.�/�)�*�&�'�#�$�!�"�(�)�'�(�%�&�$�%�#�$�!�"�)�*�&�'�"�#� �!� � �"�"�$�$�&�&�(�(�*�*�3�3�-�-�/�/�1�1�3�3�4�4�6�6�8�8�:�:�<�<�>�>�@�@�A�A�C�C�E�E���������   $               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���-���^���e����{{{����"""�'''�***�222�777�999�:::�333�777�:::�@@@�CCC�FFF�HHH�KKK�MMM�MMM�NNN�JJJ�DDD�EEE�EEE�DDD�EEE�EEE�EEE�OOO�QQQ�QQQ�RRR�RRR�RRR�NNN�NNN�NNN�NNN�NNN�PPP�JXJ�E^E�FcG�DfE�CiD�AlB�AqB�?t@�@yA�?}@�<~=�=�>�9�:�6�7�2�3�,�-�*�+�'�(�-�.�,�-�*�+�(�)�'�(�%�&�$�%�.�/�+�,�%�&�$�%�!�"�"�"�$�$�&�&�(�(�5�5����n�q�/�/�1�1�3�3�4�4�6�6�8�8�:�:�<�<�>�>�?�?�A�A�C�C�E�E���������   #               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���-���^���d����|||����###�(((�+++�444�999�;;;�<<<�444�777�<<<�AAA�DDD�GGG�JJJ�MMM�NNN�OOO�PPP�KKK�FFF�FFF�EEE�EEE�FFF�FFF�GGG�QQQ�SSS�TTT�TTT�TTT�TTT�PPP�PPP�PPP�PPP�PPP�MTM�JZJ�I]I�IbI�IfJ�FhG�FlG�FqG�CsD�CxD�D}E�@~A�A�B�>�?�<�=�7�8�0�1�/�0�2�3�1�2�0�1�-�.�+�,�)�*�(�)�'�(�3�4�0�1�(�)�&�'�"�#�"�#�$�$�&�&�2�3�����������o�r�1�1�2�2�4�4�6�6�8�8�:�:�<�<�>�>�?�?�A�A�C�C�E�E���������   !               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���-���^���d����|||����$$$�)))�,,,�666�:::�<<<�===�555�888�<<<�BBB�FFF�III�LLL�NNN�QQQ�QQQ�RRR�MMM�GGG�GGG�GGG�GGG�GGG�GGG�HHH�SSS�UUU�VVV�VVV�VVV�VVV�RRR�RRR�QQQ�RRR�RSR�PVP�NYN�N^N�NbN�MfM�JgK�IkJ�JpK�HsI�GwH�H}I�E~F�G�H�C�D�@�A�<�=�6�7�8�9�7�8�5�6�4�5�1�2�.�/�,�-�+�,�*�+�7�8�6�7�+�,�)�*�$�%�#�$�$�%�1�1�������������ئ���q�s�2�2�4�4�6�6�8�8�:�:�<�<�=�=�?�?�A�A�C�C�E�E���������               
   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���-���]���d����xxx����$$$�+++�---�777�<<<�>>>�???�666�999�>>>�CCC�GGG�III�LLL�OOO�RRR�SSS�SSS�NNN�HHH�III�HHH�III�III�III�III�VVV�WWW�WWW�YYY�XXX�WWW�SSS�SSS�TTT�TTT�TTT�STS�SYS�Q\Q�RbR�PdP�NgN�MjN�NpO�MsN�MxN�M}N�I~J�L�M�H�I�E�F�A�B�>�?�=�>�;�<�9�:�8�9�5�6�1�2�/�0�.�/�-�.�=�>�:�;�.�/�,�-�&�'�$�%�/�0��ۇ�����KpK�ݜJ���ا���r�t�4�4�6�6�8�8�:�:�;�;�=�=�?�?�A�A�C�C�D�D���������               
   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���-���]���dyyy�rrr����%%%�,,,�...�999�>>>�@@@�AAA�666�:::�???�EEE�HHH�KKK�NNN�QQQ�SSS�VVV�VVV�PPP�JJJ�JJJ�JJJ�JJJ�KKK�KKK�KKK�WWW�YYY�ZZZ�YYY�ZZZ�ZZZ�UUU�UUU�UUU�UUU�VVV�UUU�VWV�V\V�VaV�VfV�SgS�QjQ�SpT�QsR�RxS�S~T�N~O�Q�R�N�O�J�K�H�I�B�C�@�A�?�@�=�>�<�=�8�9�5�6�3�4�1�2�0�1�A�B�?�@�1�2�0�1�'�)�.�/�؄���ګ�HcH      
��F���ק���s�u�6�6�8�8�:�:�;�;�=�=�?�?�A�A�C�C�D�D���������               	   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���-���]���dsss�mmm����&&&�---�000�;;;�@@@�BBB�BBB�777�:::�???�FFF�JJJ�LLL�OOO�RRR�VVV�WWW�XXX�RRR�LLL�LLL�KKK�KKK�LLL�LLL�LLL�YYY�[[[�[[[�\\\�\\\�[[[�VVV�VVV�WWW�VVV�XXX�WWW�XXX�XYX�Z`Z�YdY�VfV�WkW�XqX�UrV�VxW�X~Y�TU�W�X�T�U�R�S�N�O�F�G�D�E�C�D�A�B�@�A�;�<�8�9�6�7�5�6�3�4�F�G�C�D�5�6�3�4�3�4�ԁ���ԫ宔@O@             ��D���ب���t�w�8�8�9�9�;�;�=�=�?�?�A�A�B�B�D�D���������                  ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���,���\���cmmm�ggg����&&&�...�111�<<<�BBB�DDD�DDD�888�<<<�AAA�FFF�KKK�NNN�PPP�SSS�WWW�ZZZ�ZZZ�TTT�LLL�MMM�LLL�LLL�MMM�MMM�NNN�[[[�]]]�]]]�^^^�^^^�^^^�YYY�XXX�YYY�YYY�YYY�XXX�ZZZ�[[[�^_^�]c]�[f[�ZjZ�[o[�ZsZ�[x\�]^�YZ�\�]�Z�[�W�X�S�T�K�L�I�J�G�H�F�G�D�E�?�@�;�<�:�;�8�9�7�8�K�L�I�J�8�9�@�A�|�~�ܝΧڪ�.B.'         	         ���D���٩���v�x�9�9�;�;�=�=�?�?�A�A�B�B�D�D���������            	      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���,���\���cfff�aaa����'''�///�222�===�DDD�EEE�EEE�999�===�AAA�HHH�LLL�OOO�QQQ�TTT�WWW�[[[�]]]�UUU�MMM�NNN�NNN�NNN�NNN�OOO�OOO�\\\�___�___�```�___�```�ZZZ�ZZZ�ZZZ�ZZZ�ZZZ�ZZZ�[[[�]]]�aaa�aba�`f`�_j_�aqa�^r^�`y`�d�e�_�`�b�c�`�a�]�^�W�X�O�P�M�N�L�M�J�K�G�H�B�C�?�@�=�>�<�=�:�;�R�S�M�N�D�E�Ѐ�۟Рͤ�&1&/                        ���C���٩���w�z�;�;�=�=�?�?�@�@�B�B�N�N���������                  ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���,���\���b___�[[[����(((�000�222�???�EEE�GGG�HHH�999�>>>�BBB�JJJ�LLL�PPP�SSS�VVV�YYY�\\\�^^^�VVV�NNN�OOO�OOO�OOO�OOO�OOO�PPP�^^^�aaa�```�bbb�aaa�aaa�\\\�\\\�\\\�]]]�]]]�\\\�\\\�^^^�ccc�eee�efe�bhb�fqf�csc�eye�i�i�d�e�h�i�f�g�c�d�]�^�S�T�R�S�P�Q�N�O�L�M�F�G�B�C�A�B�?�@�>�?�U�V�X�Y�~΀�ݩܬί�% 7   %                           ���C���٪���x�z�=�=�?�?�@�@�B�B�d�f���������         	         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���,���\���bXXX�UUU���   �)))�111�444�AAA�GGG�III�III�:::�>>>�CCC�KKK�NNN�QQQ�TTT�VVV�ZZZ�]]]�___�XXX�PPP�QQQ�PPP�OOO�PPP�PPP�PPP�```�bbb�ccc�ddd�ddd�ddd�^^^�^^^�^^^�^^^�^^^�___�^^^�```�ddd�fff�fff�ghg�jpj�iti�jzj�n�n�j�j�o�p�m�n�i�j�c�d�Y�Z�W�X�U�V�R�S�P�Q�J�K�F�G�D�E�C�D�A�B�`�a��ˆ��ק���Ży{y`   0   %                              ���C���ګ���z�|�>�>�@�@�B�B�|�~���������   
   	            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���,���[���bRRR�SSS���   �)))�111�444�BBB�III�KKK�JJJ�:::�???�DDD�KKK�OOO�RRR�UUU�XXX�[[[�___�aaa�ZZZ�QQQ�RRR�PPP�QQQ�PPP�RRR�RRR�bbb�ddd�fff�fff�fff�eee�___�___�___�___�```�___�```�aaa�eee�hhh�hhh�jjj�opo�ntn�p{p�t�t�o�o�t�t�s�t�n�o�j�k�_�`�\�]�Z�[�W�X�U�V�O�P�I�J�H�I�F�G�H�I��ǈ��Ӯ���º����qqq[   0   %                                  ���C���۫���{�}�@�@�D�D����������U                  ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���,���[���aYYY�XXX���   �***�333�555�DDD�KKK�MMM�MMM�;;;�???�DDD�LLL�PPP�SSS�VVV�YYY�\\\�___�ccc�[[[�QQQ�RRR�RRR�RRR�RRR�SSS�SSS�ddd�fff�ggg�ggg�hhh�ggg�aaa�aaa�aaa�aaa�aaa�aaa�aaa�bbb�fff�iii�iii�lll�qqq�sts�tzt�z�z�u�u�|�|�y�y�v�w�o�p�d�e�a�b�^�_�[�\�Z�[�S�T�M�N�L�M�M�N�p�q��ɨ�������������rrrZ   /   $                                      ���B���ڬ���|�~�t�v���������g�g                  ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���,���[���a___�^^^���   �+++�444�777�FFF�MMM�OOO�NNN�;;;�@@@�EEE�MMM�QQQ�TTT�XXX�ZZZ�]]]�aaa�ddd�]]]�SSS�SSS�SSS�SSS�TTT�TTT�UUU�eee�iii�jjj�iii�jjj�iii�bbb�ccc�ccc�bbb�ccc�ccc�ccc�ccc�hhh�jjj�lll�nnn�sss�uuu�{|{�����|�|�������{�{�v�w�i�j�f�g�c�d�`�a�_�`�W�X�Q�R�Q�R�m�n���������������������qqqY   /   $                     ��� ���              ���B���ۭ�������������D                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���+���Z���afff�ddd���   �+++�444�888�GGG�NNN�QQQ�PPP�<<<�@@@�GGG�NNN�RRR�UUU�YYY�[[[�^^^�bbb�eee�^^^�TTT�UUU�TTT�TTT�UUU�UUU�UUU�ggg�kkk�jjj�kkk�kkk�kkk�ddd�ddd�eee�eee�eee�ddd�fff�eee�jjj�lll�mmm�ooo�ttt�vvv����������������������}�}�n�o�k�l�i�j�e�f�d�e�Z�[�W�X�l�m�������������������������qqqY   /   $                     ��� ���                  ���B���ۨ������                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���+���Z���ammm�jjj���!!!�,,,�666�999�HHH�QQQ�QQQ�QQQ�===�@@@�GGG�OOO�RRR�VVV�YYY�]]]�```�ccc�ggg�___�UUU�UUU�VVV�TTT�UUU�UUU�VVV�iii�lll�mmm�mmm�mmm�lll�fff�eee�fff�fff�eee�fff�fff�fff�kkk�mmm�nnn�qqq�vvv�xxx�����������������������������t�t�p�q�m�n�k�l�i�j�a�b�l�m�}�~�����rsr�����������������qqqY   /   $                     ��� ��� ���                   ���B���Ġ�                           ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���+���Z���asss�ppp���!!!�---�777�:::�JJJ�RRR�TTT�SSS�>>>�BBB�HHH�PPP�SSS�WWW�ZZZ�]]]�```�ddd�hhh�```�VVV�VVV�WWW�VVV�VVV�VVV�WWW�kkk�ooo�ooo�nnn�ppp�ooo�ggg�hhh�hhh�ggg�hhh�hhh�ggg�ggg�mmm�nnn�ppp�rrr�xxx�zzz�����������������������������x�x�v�v�s�t�p�q�o�p�o�p�{�{�����uuu�sss�����������������pppY   /   $                     ��� ��� ��� ��� ���                 ��                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���+���Y���`zzz�uuu��   �!!!�---�888�;;;�LLL�TTT�WWW�UUU�>>>�AAA�GGG�QQQ�TTT�XXX�[[[�___�aaa�fff�iii�aaa�XXX�XXX�WWW�VVV�WWW�WWW�XXX�mmm�ppp�ppp�qqq�rrr�qqq�hhh�iii�iii�iii�iii�iii�jjj�iii�mmm�qqq�ppp�sss�zzz�zzz�����������������������������~�~�|�|�w�w�w�x�y�z�~�~�����uuu�ttt�ttt�����������������pppY   /   $                     ��� ��� ��� ��� ��� ��� ���                                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���+���Y���`����|||��   �"""�...�888�;;;�NNN�VVV�XXX�WWW�???�CCC�III�QQQ�UUU�YYY�\\\�___�bbb�fff�jjj�ccc�XXX�YYY�XXX�XXX�XXX�YYY�YYY�ooo�rrr�sss�sss�rrr�rrr�jjj�jjj�jjj�kkk�kkk�lll�kkk�kkk�ooo�rrr�qqq�ttt�{{{�}}}���������������������������������������|�|���������xxx�vvv�ttt�uuu�����������������pppY   /   $                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���+���Y���_����|||��!!!�###�///�:::�<<<�PPP�YYY�ZZZ�XXX�???�CCC�HHH�RRR�VVV�YYY�\\\�```�ddd�ggg�kkk�aaa�YYY�ZZZ�XXX�YYY�YYY�YYY�ZZZ�ppp�sss�ttt�ttt�vvv�ttt�kkk�lll�lll�mmm�lll�mmm�mmm�mmm�qqq�rrr�ttt�uuu�|||�~~~�����������������������������������������������������www�www�vvv�vvv�����������������pppY   /   $                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���+���X���_����}}}��!!!�###�///�;;;�>>>�QQQ�ZZZ�\\\�ZZZ�>>>�CCC�III�SSS�WWW�[[[�^^^�```�ddd�iii�kkk�ccc�ZZZ�[[[�ZZZ�YYY�[[[�[[[�ZZZ�qqq�uuu�vvv�vvv�www�vvv�nnn�mmm�mmm�nnn�nnn�nnn�mmm�mmm�rrr�uuu�ttt�www�~~~���������������������������������������������������������xxx�xxx�www�www�zzz�|||���������oooY   /   $                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���*���X���_����}}}��"""�###�000�;;;�>>>�RRR�\\\�^^^�\\\�???�CCC�JJJ�SSS�XXX�[[[�___�bbb�eee�iii�mmm�ddd�ZZZ�\\\�[[[�YYY�ZZZ�[[[�[[[�ttt�vvv�xxx�xxx�xxx�xxx�nnn�nnn�ooo�ooo�ppp�ppp�ooo�ooo�uuu�vvv�uuu�xxx�������������������������������������������������������������zzz�yyy�www�xxx�sss�uuu���������oooY   /   $                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���*���W���^����}}}��!!!�$$$�111�===�@@@�TTT�___�```�]]]�???�CCC�JJJ�TTT�XXX�\\\�___�ccc�fff�jjj�nnn�ddd�ZZZ�\\\�[[[�\\\�[[[�\\\�]]]�ttt�zzz�zzz�yyy�zzz�{{{�ppp�ooo�ooo�ppp�qqq�qqq�qqq�qqq�vvv�www�www�zzz�������������������������������������������������������������zzz�zzz�xxx�xxx�ttt�nnn���������oooY   /   $                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���*���W���^����}}}�   �"""�$$$�222�>>>�AAA�VVV�aaa�bbb�```�@@@�DDD�JJJ�UUU�YYY�]]]�___�ccc�ggg�kkk�ooo�ddd�ZZZ�]]]�\\\�[[[�\\\�\\\�]]]�vvv�{{{�{{{�{{{�{{{�{{{�qqq�qqq�rrr�rrr�rrr�sss�sss�sss�yyy�yyy�xxx�{{{�������������������������������������������������������������zzz�zzz�zzz�zzz�{{{�uuu���������oooY   /   $                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���*���W���^����}}}�   �"""�$$$�333�???�BBB�WWW�bbb�eee�bbb�@@@�DDD�KKK�UUU�ZZZ�]]]�```�eee�hhh�kkk�ooo�eee�ZZZ�]]]�]]]�\\\�]]]�\\\�]]]�www�|||�|||�}}}�}}}�~~~�sss�sss�sss�ttt�ttt�uuu�ttt�ttt�zzz�{{{�zzz�}}}�������������������������������������������������������������{{{�|||�zzz�{{{�����}}}���������oooY   /   $                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���)���W���^����}}}�   �"""�%%%�333�@@@�CCC�XXX�eee�ggg�ccc�AAA�EEE�KKK�VVV�[[[�___�aaa�eee�iii�mmm�ooo�eee�ZZZ�]]]�]]]�^^^�]]]�^^^�^^^�yyy�~~~�~~~�������ttt�uuu�ttt�uuu�uuu�uuu�ttt�vvv�zzz�|||�{{{�~~~�������������������������������������������������������������}}}�|||�{{{�{{{�����������������oooW   /   $                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���)���V���\����}}}�!!!�"""�$$$�555�BBB�DDD�[[[�hhh�iii�ddd�AAA�DDD�KKK�VVV�ZZZ�___�aaa�eee�iii�mmm�ppp�ggg�YYY�]]]�^^^�]]]�]]]�___�___�{{{������������������vvv�vvv�vvv�www�vvv�www�vvv�www�|||�~~~�|||�����������������������������������������������������������������}}}�}}}�}}}�{{{�����������������oooW   .   #                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���)���U���\����}}}�!!!�###�%%%�555�CCC�EEE�\\\�hhh�kkk�fff�AAA�EEE�LLL�WWW�\\\�___�bbb�fff�jjj�nnn�qqq�fff�YYY�]]]�^^^�^^^�^^^�___�aaa�}}}���������������������vvv�www�vvv�www�www�www�xxx�xxx������}}}�����������������������������������������������������������������~~~�}}}�|||�|||�����������������oooV   -   "                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 ���(���T���Z����}}}�"""�$$$�%%%�666�DDD�FFF�^^^�kkk�nnn�hhh�@@@�EEE�LLL�XXX�]]]�___�ccc�fff�kkk�nnn�rrr�fff�ZZZ�\\\�^^^�___�```�```�```�~~~���������������������xxx�yyy�xxx�xxx�yyy�zzz�zzz�zzz���������������������������������������������������������������������������~~~�~~~�~~~�����������������qqqT   ,   !         
            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 ���'���S���Y����~~~�###�$$$�%%%�777�EEE�GGG�___�nnn�ppp�jjj�@@@�DDD�LLL�YYY�]]]�```�ddd�ggg�kkk�nnn�sss�fff�YYY�^^^�^^^�___�aaa�```�aaa����������������������zzz�zzz�zzz�{{{�zzz�zzz�{{{�zzz�������������������������������������������������������������������������������~~~�}}}�����������������uuuR   )            	             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 ���'���R���X����}}}�###�%%%�&&&�888�FFF�III�aaa�ppp�rrr�mmm�@@@�FFF�MMM�XXX�^^^�aaa�ddd�hhh�lll�ppp�sss�fff�ZZZ�]]]�^^^�___�```�```�bbb�������������������������{{{�|||�{{{�|||�|||�|||�|||�|||������������������������������������������������������������������������������~~~�~~~�}}}�����������������yyyO   &            	             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                         ��� ��� ��� ��� ��� ���                 ���%���P���U����~~~�$$$�&&&�&&&�888�HHH�KKK�ccc�sss�ttt�ooo�AAA�FFF�MMM�YYY�^^^�aaa�ddd�hhh�lll�qqq�sss�ggg�YYY�]]]�^^^�```�aaa�bbb�bbb�������������������������|||�}}}�}}}�}}}�}}}�}}}�}}}�~~~�����������������������������������������������������������������������������~~~�}}}�|||�{{{��������������������K   #                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                 ��� ��� ��� ���                  ���$���N���S����~~~�$$$�&&&�'''�999�JJJ�LLL�ddd�ttt�vvv�qqq�AAA�EEE�NNN�ZZZ�^^^�bbb�eee�iii�mmm�ppp�uuu�ggg�YYY�^^^�^^^�___�aaa�bbb�bbb�������������������������}}}�}}}�~~~�~~~�~~~�����������������������������������������������������������������������������������}}}�{{{�{{{�{{{�������������������F            
                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                          ��� ���                  ���"���L���P��������&&&�'''�(((�:::�KKK�NNN�ggg�www�yyy�rrr�AAA�FFF�MMM�[[[�___�bbb�fff�jjj�nnn�qqq�vvv�iii�YYY�]]]�^^^�```�aaa�ccc�ccc����������������������������������������������������������������������������������������������������������������������������}}}�{{{�{{{�zzz���������������z���A            	                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                          ��� ���              ���!���J���N��������CCC�'''�(((�<<<�LLL�OOO�iii�yyy�|||�ttt�AAA�FFF�MMM�ZZZ�___�bbb�fff�jjj�ooo�rrr�uuu�iii�XXX�\\\�]]]�___�bbb�ddd�ccc����������������������������������������������������������������������������������������������������������������������������������{{{�zzz�yyy����������������y���v���;         
                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                             ������H���L���ć���uuu�AAA�***�===�NNN�PPP�jjj�|||�~~~�www�AAA�EEE�NNN�[[[�```�ccc�ggg�kkk�nnn�rrr�xxx�iii�YYY�]]]�]]]�___�bbb�ccc�ddd�������������������������������������������������������������������������������������������������������������������������������������zzz�zzz��������������������t���q���.                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                            ������H���J���N������������������������������������������������������������������������������������������������������������������������������������������������������ttt�iii�eee�ppp�|||����������������������������������������������������������������������������������������������������s���o���mddd                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                      	   
      
   	                                            ���-���H���K���O���ǌ��򋋋���������������������������������������������������������������������������������������������������������������������������������������������vvv�iii�]]]�ggg�ttt������������������������������������������������������������������������������������������������r���n���k���F   
                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                	                        
                                    iii���5���J���M���O���T���[����а�׿�����鉉�������������������������������������������������ٝ��|���u���o���i���e���a���^���]���\���\���[���[���\���\���]���]���^���^���^���_���_���`���b���c���g���k�����������������������������������������������������������������������z���u���p���m���j���L\\\                          ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                  ������/���;¿�D���r�ͦ�ڷ|�ɥg}����{{{�����������������������������������������}}}�����i���a���Y���R���L���G���D���A���@���?���@���@���@���@���@���A���A���A���A���B���B���D���E���G���K���O�����������������������������������������������������������v���o���g���`���Y���R���B���(   	                          ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���             
���+�γ�F<2                           	                                 	      OD9�ĬW翄�י:s�v _�qbqme�\\\�������������������������������������kkk�\\\�___�   A   6   +   !               	                                          	         bbb�\\\�������������������������������������___�\\\�999|   H   =   2   '            
                          ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���          	   �д��Ѱ��̰�7/'                            	                           	   
   SSG�ȳ^�Ŋ��=z�} d�v d�tfrmd�\\\�������������������������������������kkk�\\\�``^�   @   5   *                                                                	      bbb�\\\�������������������������������������___�\\\�999|   G   <   1   %                                    ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���          	�¦d�Ҳ������ά��Ȯ�0)"%                            	                     	      [OO�̴h�Ǝ��?�Ձ k�| i�x h�sksmd�\\\�������������������������������������kkk�\\\�a`^� C   4   )                                                                     bbb�\\\�������������������������������������___�\\\�999{   F   ;   0   $                             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       �� �ѳ��Ě��v���d��ϭ��Ǭ�*$*   #   !                        	         	   
      ^SI�Ͷp�Ǒ��A�ۂ r� o�} n�x m�vosmc�\\\�������������������������������������kkk�\\\�ca]�! F 8   )            
                                                           bbb�\\\�������������������������������������___�\\\�999{   F   ;   /   $                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       �ǫv�ѳ���7��q ��r ���e��έ��ū�("-   %   #                                    aWM�εx�Ȕ��C�߁ zۂ x� t�z s�x r�vtsmc�\\\�������������������������������������kkk�\\\�db]�1# J' ; .                                              ��� ���                       bbb�\\\�������������������������������������___�\\\�999{   F   ;   /   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       	�̮��ѱ��r��p ��q ��q ���d��Ϭ��é�&!/   '   #                               `OF�͵��ɖ��C�� ��� �� |� {�{ x�v v�wytmc�\\\�������������������������������������kkk�\\\�ec\�>* N8( @. 2# $                                       ��� ��� ���                       bbb�\\\�������������������������������������___�\\\�999{   F   ;   /   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       	�ή������n ��o ��p ��p ��q ���c��Ϭ�����%1   (   $   !                     ZRJ�δ��ș��F�� �� ��� �� ��| �| }�w |�u}unb�\\\�������������������������������������kkk�\\\�gc\�H2 QG1 DB/ 6:& (-$                                         ��� ���                       bbb�\\\�������������������������������������___�\\\�999{   F   ;   /   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �|c�а���n��m ��m ��o ��o ��p ��p ���c��ϭ��¨�$2   (   %   !               UN@$�˳��ʜ��F�� ��~ �� ��} ��~ ��} ��z ��y ��w�unb�\\\�������������������������������������kkk�\\\�hd\�S8 VQ9 HR8 ;O8 -G0  ;/                                     ��� ���                       bbb�\\\�������������������������������������___�\\\�999{   F   ;   /   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ͦ�(�ͮ���Y��l ��l ��m ��n ��o ��p ��p ���c��ή�����$2   )   &   #   !      RE?)�̲��ɞ��G��} ��} ��} ��} ��~ ��| ��| ��{ ��w ��y�vnb�\\\�������������������������������������kkk�\\\�hd[�^? Z^@ L^B >bC 2aF %Z< L= FFF+++                           ��� ���                       bbb�\\\�������������������������������������___�\\\�999{   F   ;   /   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    Ȝ�)�̬���W��k ��k ��l ��m ��n ��o ��o ��p ���c��Ϯ�����#3   *   (   %   #MB7.�ɱ��ʠ��H��{ ��{ ��| ��| ��| ��| ��} ��{ ��z ��y ��w�vna�\\\�������������������������������������kkk�\\\�je[�fE ]iF PlI BoM 5sO *wU pJ ��[���                            ��� ���                       bbb�\\\�������������������������������������___�\\\�999{   F   ;   /   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    Ȝ�)�˪���V��i ��k ��k ��l ��m ��n ��o ��o ��p ���b��έ��§�#4   ,   *E;64�ȭ��ʢ���I��z ��z ��z ��z ��{ ��{ ��{ ��{ ��{ ��y ��x ��y�wna�\\\�������������������������������������kkk�\\\�ke[�oJ `qM SwP F|T 9�Y .�_ #�k
īr���                        ��� ��� ���                       bbb�\\\�������������������������������������___�\\\�999{   F   ;   /   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    Ȝ�)�ʩ���U��h ��i ��j ��k ��l ��l ��n ��n ��o ��p ���b��Ϯ�����"5B90:�Ƭ��ͥ���J��x ��y ��y ��y ��z ��z ��{ ��{ ��z ��z ��z ��w ��y�xna�\\\�������������������������������������kkk�\\\�mfY�vM c{R W�V J�[ >�b 1�j &Ȣ\/Ҽ�#��u                        ��� ��� ���                       bbb�\\\�������������������������������������___�\\\�999{   F   ;   /   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    Ȝ�)�ȧ���T��g ��h ��i ��j ��k ��l ��l ��n ��n ��o ��p ���b��ϯ��¨��Ƭ��ͩ���K��v ��v ��x ��x ��y ��y ��y ��y ��z ��z ��z ��y ��x ��w�xn`�\\\�������������������������������������kkk�\\\�nfY�~R g�U Z�[ O�b A�h 6ȤX@Ѻ�7���                                                           bbb�\\\�������������������������������������___�\\\�:::{   F   :   /   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ę{*�ǥ���S��f ��g ��h ��i ��j ��k ��l ��l ��n ��n ��o ��p ���b��Я��Ϋ���K��s ��u ��u ��u ��w ��x ��y ��y ��y ��y ��z ��y ��x ��w ��y�yn`�\\\�������������������������������������kkk�\\\�ngYՅU l�Y _�] R�e FŠSSҶ�I���$                                                         bbb�\\\�������������������������������������___�\\\�:::{   F   :   /   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ę{*�ţ���S��f ��f ��g ��h ��i ��j ��k ��k ��l ��n ��n ��o ��p ���b���M��r ��s ��s ��u ��u ��u ��w ��w ��x ��y ��x ��x ��y ��x ��w ��{�zo_�\\\�������������������������������������kkk�\\\�pgX֊W o�\ d�a WRf̳�\���1      	                                                	      bbb�\\\�������������������������������������___�\\\�:::{   E   :   .   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ē{*�ġ���R��e ��f ��f ��g ��h ��i ��j ��k ��k ��l ��n ��n ��o ��p ��p ��r ��r ��s ��s ��u ��u ��u ��w ��w ��x ��x ��x ��x ��x ��z��z
�zo_�\\\�������������������������������������kkk�\\\�qhX؏Z t�^h��Ryɰ�p���?                                                      	         bbb�\\\�������������������������������������___�\\\�:::{   D   9   -   "         
             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ē{*�à���Q��d ��e ��f ��f ��g ��h ��i ��j ��k ��k ��l ��m ��n ��o ��p ��p ��q ��r ��s ��s ��u ��u ��u ��w ��w ��x ��x ��x ��{��{��z	�{o_�\\\�������������������������������������kkk�\\\�rhWڕ^z��Q�Ū�����N                	                                 	   
            bbb�\\\�������������������������������������___�\\\�:::z   D   8   ,   !         
             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ē{*������P��c ��d ��e ��f ��f ��g ��h ��i ��j ��k ��k ��l ��m ��n ��o ��p ��p ��q ��r ��s ��s ��u ��u ��u ��w ��w ��x ��{��z��z��z	�{n_�\\\�������������������������������������mmm�]]]�tiW���Q�è����y_,   #                                                                bbb�\\\�������������������������������������___�\\\�;;;y   B   7   +   !         	             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��r*������O��b ��c ��d ��e ��f ��f ��g ��h ��i ��j ��k ��k ��l ��m ��n ��o ��p ��p ��q ��r ��s ��s ��u ��u ��u ��w ��{��|��z��z��y�{o_�]]]�������������������������������������ppp�```��wi�ĩ���~so:   1   )   "                                                         !   'aaa�\\\�������������������������������������___�\\\�;;;w   A   6   *            	             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��r*������N��a ��b ��c ��d ��e ��f ��f ��g ��h ��i ��j ��k ��k ��l ��m ��n ��o ��p ��p ��q ��r ��s ��s ��u ��u��y��{	��{��z��z��z��q]�___�������������������������������������yyy�ccc�}xsw�K   ?   7   0   *   %   "                                             !   $   )   /```�\\\�������������������������������������]]]�\\\�%%%a   ?   3   (            	             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��r*�����M��` ��a ��b ��c ��d ��e ��f ��f ��g ��h ��i ��j ��k ��k ��l ��m ��n ��o ��p ��p ��q ��r ��s ��s��y	��z
��y	��{��y��z��{��wV�bbb�|||�������������������������������������fff�onn�!!!\SI@   9   3   /   ,   )   (   '   &   &   &   &   &   &   &   &   '   (   )   +   .   2   7]]]�\\\�������������������������������������\\\�]]]�   G   <   1   &                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��r*�����L��` ��` ��a ��b ��c ��d ��e ��f ��f ��g ��h ��i ��j ��k ��k ��l ��m ��n ��o ��p ��p ��q ��r��x
��z��z
��z	��y��y��{	��}��~L�ddd�sss�������������������������������������hhh�iii�>>>x"""[SK   B   =   9   6   4   3   2   1   1   1   1   1   1   1   1   2   3   4   6   9   =]]]�\\\�```�������������������������������������\\\�^^^�   D   9   .   #                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��l*������K��_ ��` ��` ��a ��b ��c ��d ��e ��f ��f ��g ��h ��i ��j ��k ��k ��l ��m ��n ��o ��p ��r��v��x��z��x
��z	��y��z
��~���̓3�fff�kkk�������������������������������������vvv�iii�mmm�'''b!!!\UN   G   D   A   @   ?   >   =   =   =   =   =   =   =   =   >   >   ?   A   D111e___�\\\�}}}�������������������������������������\\\�___�   @   6   *             
            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��l*�����K��^ ��_ ��` ��` ��a ��b ��c ��d ��e ��f ��f ��g ��h ��i ��j ��k ��k ��l ��m ��n ��p��v
��x��x��x��x
��x	��z	��|��~�����nnm�kkk�����������������������������������������mmm�jjj�mmm�XXX�]XQ   M   L   J   I   H   H   H   H   H   H   H   H   H   H   I   JS\\\�^^^�\\\�fff�������������������������������������nnn�\\\�aaa�   <   1   '            	             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��l*�����J��] ��^ ��_ ��` ��` ��a ��b ��c ��d ��e ��f ��f ��g ��h ��i ��j ��k ��k ��l ��o��u��v��w��w��x��w
��x��y��~������ Ƅyn�mmm���������������������������������������������ppp�iii�hhh�fff�fff�ccc�___�```�```�```�```�```�```�```�```�```�```�```�```�```�```�___�]]]�\\\�\\\�hhh�����������������������������������������___�\\\�SSS�   7   ,   #                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��j+�����I��\ ��] ��^ ��_ ��` ��` ��a ��b ��c ��d ��e ��f ��f ��g ��h ��i ��j ��k ��l��s��v��v��v��v��w
��v	��w
��z��}������ȵ�Y�ooo�vvv����������������������������������������������mmm�fff�ddd�```�]]]�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�ddd����������������������������������������������\\\�^^^�   ;   1   (            
                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��j+�����H��[ ��\ ��] ��^ ��_ ��` ��` ��a ��b ��c ��d ��e ��f ��f ��g ��h ��i ��k��r��s��t��u��v��u��v
��u
��x��z��~������!��*�xvt�sss�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ddd�\\\�bbb�   5   ,   "                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��d+�����G��Z ��[ ��\ ��] ��^ ��_ ��` ��` ��a ��b ��c ��d ��e ��f ��f ��g ��i��p��s��s��s��s��u��u��u��u
��x��z��~�������$��+ΰ�d�ttt�~~~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������\\\�^^^�E   /   %            
                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��d+�����F��Y ��Z ��[ ��\ ��] ��^ ��_ ��` ��` ��a ��b ��c ��d ��e ��f ��g��o��q��r��r��s��r��s��t��u��t
��w��z��~�������%���*��4Ђ�~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������```�\\\�aaa�   0   (                               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��d+�����E��Y ��Y ��Z ��[ ��\ ��] ��^ ��_ ��` ��` ��a ��b ��c ��d ��f��n��p��p��q��q��r��r��r��r��t��s
��v��z��}���� ��%��,�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ddd�\\\�```�4   )   !            	                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��d+�����D��X ��Y ��Y ��Z ��[ ��\ ��] ��^ ��_ ��` ��` ��a ��b ��d��m��p��p��p��p��p��q��q��r��q��r��s
��u��y��|���� ��'������׽��ʷ�������������������������������������������������������������������������������������������������������������������������������������������������������������������������iii�\\\�___�000K   )   !            
                    ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��d+�����D��W ��X ��Y ��Y ��Z ��[ ��\ ��] ��^ ��_ ��` ��` ��b��l��n��o��o��p��o��p��p��q��q��r��q
��r
��u��x��{�����������׽��ȳ���X���e���ݘ�����������������������������������������������������������������������������������������������������������������������������������������������������������ccc�\\\�^^^�TTTs   (   !                               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��^+�����C��V ��W ��X ��Y ��Y ��Z ��[ ��\ ��] ��^ ��_ ��a��j��m��n��n��n��o��o��o��o��p��p��q��q
��q	��s��x��y��}������y��׾��͵˄}X���]���k���Ӗ�����������������������������������������������������������������������������������������������������������������������������������������������|||�___�\\\�___�QQQm   %                                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �~`*�����B��U ��V ��W ��X ��Y ��Y ��Z ��[ ��\ ��] ��_��j��m��l��m��m��n��n��n��o��n��o��o��p��p
��q
��q��u��x��{��~��� ���z��ٿ��̷͉��Y���_���h��������������������������������������������������������������������������������������������������������������������������������������������ccc�\\\�\\\�```�555C   "                                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �~`*�����A��T ��U ��V ��W ��X ��Y ��Y ��Z ��[ ��]��i��l��l��l��l��l��m��m��n��n��n��n��n��o��o
��p
��q
��s��v��z��|�����"���|��ٿ��η̇��X���Y���^���z����zzz�uuu�sss�zzz�������������������������������������������������������������������������������������������������}}}�lll�]]]�\\\�\\\�^^^�ddd�%                  
                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    āb*��~��@��S ��T ��U ��V ��W ��X ��Y ��Y ��[��g��k��k��k��l��l��k��l��l��m��m��n��n��m��n��n��o
��o	��r��t��w��z��}�����!���{��ؾ��η̇�U}}}P���O���O���|||�sss�ooo�mmm�jjj�hhh�eee�ccc�```�]]]�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�___�eee�###*                     	                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ͆`(��|��~?��S ��S ��T ��U ��V ��W ��X ��Z��f��i��j��j��j��k��k��l��k��k��l��l��m��m��m��m��m��n
��n	��p
��r��v��w��{��~������ ���{��ؽ��ͷ́||QyyyJ{{{H|||F~~~D���H����xxx�qqq�kkk�ggg�aaa�___�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�]]]�^^^�```�aaa�eee�YYYc                        	                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �sS��z��F��R ��S ��S ��T ��U ��V ��X��e��i��i��i��i��j��j��j��k��k��k��k��k��l��l��m��m��m��m
��m	��n��p
��s��v��w��z��}��������x��׽��ε�}wwLpppBppp@sss<uuu9rrr5rrr1sss.ppp*ggg']]]-ZZZ4WWW3ZZZ4ZZZ4ZZZ4ZZZ4WWW3WWW3SSS2PPP1III/AAA.<<<-888,888,888,                                 	                             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ��w��]��Q ��R ��S ��S ��T ��V��d��h��h��i��h��h��i��i��i��j��j��k��j��k��k��k��l��l��m��l
��m	��m��n��p��s��v��v��z��}��~�����x��ֺ��̵�yrrDiii:hhh6jjj2hhh,ggg'ddd$ZZZFFF...                                          	                                   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ��v���s��Q��Q ��R ��S ��T��c��g��g��g��h��h��h��h��h��i��i��i��j��j��j��j��j��k��k��l��l
��l
��l	��m��n��p
��r��u��w��y��z��}��}���v��չ��Ͳ�skk;^^^1bbb,]]]']]]!TTTGGG---            
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   	   	   	                                             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ��r���v��^��P ��Q ��S��c��f��f��f��g��g��g��h��g��g��h��h��i��i��i��j��i��j��j��j��k��k
��l
��k	��l��l��n��o	��r
��s��v��w��y��y��{���s��Է��˱�pff1QQQ&OOO MMM>>>000      	                                                                                                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       �j<��u��R��O ��Q��a��e��f��e��f��f��f��g��g��g��g��g��g��h��h��h��i��i��i��i��j��j��j��k
��k	��k��k��l��l��n��o��r	��s��v��v��x��x���p��ӵ��̰�ic\&<<<444"""                                                                                                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���          ��r���t��m,��`��d��e��e��e��e��e��e��f��f��f��g��f��g��g��g��h��h��h��i��h��i��i��j��j
��j	��k��j��k��k��l��n��n��o��q��s��t��u��v���o��Ҵ��̯�`WN                                                                                                       ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���          �gE��q���x��l*��d��d��d��e��e��d��e��e��e��f��f��f��f��f��f��g��g��h��h��h��h��h��i��i
��j	��j��j��j��j��k��k��m��m��n��n��p��q��s��s���j��Ѳ��ͮ�m`R   	                                                                                                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���              �i=��s���|�فG��c��c��d��d��d��d��d��d��e��e��e��f��e��f��f��f��g��g��g��h��g��h��h
��i	��i��j��j��j��j��j��k��l��m��m��n ��o ��q ��r �����ɤ��в��ͯ�                          ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 �k4��p���}��i��v8��g#��c��c��d��c��d��d��d��e��e��e��e��e��f��f��f��g��g��g��g��g
��h	��h	��i��i��j��i��j��j��j��l��l��m ��n��~���X��˩��έ��ʬ��zk                       ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 �^F��p���w����������x��c��^��_��^��_��`��`��_��`��`��a��a��a��b���b���b���c���c���d���c���d���d���d���e���e���f���f���g���g���i�����Ġ��ɨ��ʪ��ʨ�巜8                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                     �f*��og��r���w���x���{���|���~�����������������������������������������������������������������������������������������������à��Ţ��š��ģ��¡��M`@@                             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                                                                                                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��������������������������������������������������������������������������������������������������������������������������    �����������    �����������    �����������    �����������     �����������     ����������     ����������     ?����������     ?����������     ?�����������    ?�����������    ?�����������    ?�����������    ?�����������    ?�����������    ?�����������    ?�����������    ?�����������    ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����         ` ?����         � ?����        � ?����        � ?����        � ?����        � ?����        ��?����        ������        ������        �������        �������        �������        �������        �������        �������        �������        �������        �������        �������        �������        �������        �������        �������        �������        �������        �������        �������        �������        ?�������        �������        �������        �������        ��������       ��������� ��� ��������  ��� ��������� ��� ���������� ��� ���������� ��� ��������� ��� ������?��� ��� ��������� ��� �������� ��� �������   ��� �������   ��� �������   ��� ������ �   ��� ������ `   ��� ������     ��� ������     ��� ������     ��� ������     ��� ������     O��� ������     ��� ������     ?��� ������     ?��� ������     ��� ������     ��� ������     ?��� ������     ��  ������          ������         ������         ������         ������         ������         ������         ������        ������   �    ?������   �    ������    �    �������    |   �������    ?   �������    �����������    �����������    �����������    �����������    �����������     �����������     ����������     ?����������     ����������    ������������   ��������������������������Transparent	  TLabelLabel3LeftHTop/WidthWHeightAnchorsakLeftakBottom CaptionCopyright f�r vissa delar:  TLabelRegistrationLabelLeftHTop� Width~HeightAnchorsakLeftakBottom CaptionThis product is licensed to:  TStaticTextHomepageLabelLeftHTopHWidth� HeightCaptionhttp://XXXXXXwinscp.net/TabOrderTabStop	  TStaticTextForumUrlLabelLeftHToptWidth� HeightCaptionhttp://XXXXwinscp.net/forum/TabOrderTabStop	  TStaticTextTranslatorUrlLabelLeftHTop� Width� HeightCaptionhttp://XXXXwinscp.net/forum/TabOrderTabStop	  
TScrollBoxThirdPartyBoxLeftHTopAWidth2HeightyHorzScrollBar.Range!HorzScrollBar.VisibleVertScrollBar.Range�VertScrollBar.Smooth	VertScrollBar.Tracking	AnchorsakLeftakRightakBottom 
AutoScrollTabOrder
DesignSizeu  TLabelLabel7LeftTopWidthHeight)AnchorsakLeftakTopakRight AutoSizeCaptionTLicensavtalen f�r f�ljande program (bibliotek) �r del av applikationens licensavtal.WordWrap	  TLabelLabel4LeftTopWidth HeightCaptionLabel4Visible  TLabelPuttyVersionLabelLeftTop0Width� HeightCaption#SSH and SCP code based on PuTTY xxx  TLabelPuttyCopyrightLabelLeftTop@Width� HeightCaptionCopyright � xxx Simon Tatham  TLabelLabel8LeftTopmWidth� HeightCaption'Filemanager Toolset library Version 2.6  TLabelLabel10LeftTop}Width� HeightCaptionCopyright � 1999 Ingo Eckel  TLabelLabel1LeftTop� WidthuHeightCaptionToolbar2000 library 2.1.6  TLabelLabel2LeftTopWidth� HeightCaption$Copyright � 1998-2005 Jordan Russell  TLabelLabel5LeftTop5WidthEHeightCaptionTBX library 2.1  TLabelLabel6LeftTopEWidth� HeightCaption%Copyright � 2001-2005 Alex A. Denisov  TLabelFileZillaVersionLabelLeftTop� Width� HeightCaptionFTP code based on Filezilla xxx  TLabelFileZillaCopyrightLabelLeftTop� Width~HeightCaptionCopyright � xxx Tim Kosse  TLabelOpenSSLVersionLabelLeftTop� WidthHeightAutoSizeCaptioncThis product includes software developed by the OpenSSL Project for use in the OpenSSL Toolkit xxx.WordWrap	  TLabelOpenSSLCopyrightLabelLeftTop� Width� HeightCaption$Copyright � xxxx The OpenSSL Project  TStaticTextPuttyLicenseLabelTagLeftTopPWidthJHeightCaptionVisa licensTabOrder TabStop	OnClickDisplayLicense  TStaticTextPuttyHomepageLabelLeftTop`WidthHeightCaption5http://XXXwww.chiark.greenend.org.uk/~sgtatham/putty/TabOrderTabStop	  TStaticTextToolbar2000HomepageLabelLeftTopWidth� HeightCaption$http://www.jrsoftware.org/tb2kdl.phpTabOrderTabStop	  TStaticTextTBXHomepageLabelLeftTopUWidthzHeightCaptionhttp://www.g32.org/tbx/TabOrderTabStop	  TStaticTextFileZillaHomepageLabelLeftTop� Width� HeightCaption$http://XXXfilezilla.sourceforge.net/TabOrderTabStop	  TStaticTextOpenSSLHomepageLabelLeftTop� WidthvHeightCaptionhttp://XXX.openssl.org/TabOrderTabStop	   TButtonOKButtonLeft� Top�WidthKHeightAnchorsakRightakBottom Cancel	CaptionOKDefault	ModalResultTabOrder   TButtonLicenseButtonLeftHTop�WidthKHeightAnchorsakLeftakBottom Caption
&Licens...TabOrderOnClickLicenseButtonClick  TButton
HelpButtonLeft/Top�WidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrderOnClickHelpButtonClick  
TScrollBoxRegistrationBoxLeftHTop� Width2HeightYHorzScrollBar.VisibleVertScrollBar.Smooth	VertScrollBar.Tracking	AnchorsakLeftakRightakBottom TabOrder
DesignSize.U  TLabelRegistrationSubjectLabelLeftTopWidth!HeightAAnchorsakLeftakTopakRight AutoSizeCaptionSomeone
Somewhere, some cityWordWrap	  TLabelRegistrationLicensesLabelLeftTop+WidthkHeightCaptionNumber of Licenses: X  TStaticTextRegistrationProductIdLabelLeftTopAWidth� HeightCaptionProduct ID: xxxx-xxxx-xxxxxTabOrder OnClickRegistrationProductIdLabelClick      TPF0TAuthenticateFormAuthenticateFormLeft0TopqHelpType	htKeywordHelpKeywordui_authenticateBorderIconsbiSystemMenu BorderStylebsDialogCaptionAuthenticateFormClientHeight<ClientWidthwColor	clBtnFaceConstraints.MinHeight� Constraints.MinWidthFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameMS Sans Serif
Font.Style OldCreateOrderPositionpoMainFormCenterOnShowFormShowPixelsPerInch`
TextHeight 	TListViewLogViewLeft Top WidthwHeightAlignalClientColumnsWidth�	WidthType�   
Items.Data
.   .          ��������        Authneticating...ReadOnly		RowSelect	ShowColumnHeadersTabOrder 	ViewStylevsReport  TPanelPasswordPanelLeft TopWidthwHeight� AlignalBottomAutoSize	
BevelOuterbvNoneTabOrderVisible TPanelPromptEditPanelLeft Top WidthwHeight� AlignalTop
BevelOuterbvNoneTabOrder 
DesignSizew�   TLabelInstructionsLabelLeftTopWidthhHeight'AnchorsakLeftakTopakRight AutoSizeCaption�Instructions for authentication. Please fill in your credentials carefully. Enter all required information, including your session username and session password.XFocusControlPromptEdit1WordWrap	  TLabelPromptLabel1LeftTop8WidthhHeightAnchorsakLeftakTopakRight AutoSizeCaption&UsernameX:FocusControlPromptEdit1WordWrap	  TLabelPromptLabel2LeftTopeWidthhHeightAnchorsakLeftakTopakRight AutoSizeCaption&PasswordX:FocusControlPromptEdit2WordWrap	  TPasswordEditPromptEdit1LeftTopIWidthiHeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder   TPasswordEditPromptEdit2LeftTopvWidthiHeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder   TPanelSavePasswordPanelLeft Top� WidthwHeightAlignalTop
BevelOuterbvNoneTabOrder 	TCheckBoxSavePasswordCheckLeftTopWidthHeightCaption&�ndra l�senord till det h�rChecked	State	cbCheckedTabOrder    TPanelButtonsPanelLeft Top� WidthwHeight,AlignalTop
BevelOuterbvNoneTabOrder
DesignSizew,  TButtonPasswordOKButtonLeftvTopWidthKHeightAnchorsakTopakRight CaptionOKModalResultTabOrder   TButtonPasswordCancelButtonLeft� TopWidthKHeightAnchorsakTopakRight CaptionAvbrytModalResultTabOrder  TButtonPasswordHelpButtonLeft&TopWidthKHeightAnchorsakTopakRight Caption&Hj�lpTabOrderOnClickHelpButtonClick    TPanelBannerPanelLeft Top� WidthwHeightRAlignalBottom
BevelOuterbvNoneTabOrderVisible
DesignSizewR  TMemo
BannerMemoLeftTopWidthhHeight"AnchorsakLeftakTopakRightakBottom Color	clBtnFaceReadOnly	
ScrollBars
ssVerticalTabOrder WantReturns  	TCheckBoxNeverShowAgainCheckLeftTop5Width� HeightAnchorsakLeftakRightakBottom Caption%&Visa aldrig det h�r meddelandet igenTabOrder  TButtonBannerCloseButtonLeft� Top/WidthKHeightAnchorsakRightakBottom CaptionForts�ttModalResultTabOrder  TButtonBannerHelpButtonLeft$Top/WidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrderOnClickHelpButtonClick     TPF0TCleanupDialogCleanupDialogLeftdTop� HelpType	htKeywordHelpKeyword
ui_cleanupBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionRensa applikationsdataClientHeight+ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrder	PositionpoMainFormCenterOnShowFormShow
DesignSize�+ PixelsPerInch`
TextHeight TLabelLabel1LeftTopWidth�HeightaAnchorsakLeftakTopakRight AutoSizeCaption-  F�ljande lista inneh�ller all data som det h�r programmet lagrar p� den h�r datorn. V�lj det som du vill ska tas bort.

Om ytterligare instanser av programmet �r ig�ng, var god avsluta dem innan nedanst�ende data tas bort.

Notera att en del av dessa data kommer att �terskapas vid n�sta uppstart.WordWrap	  TButtonOKButtonLeft� TopWidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeftITopWidthKHeightAnchorsakRightakBottom Cancel	CaptionSt�ngModalResultTabOrder  	TListViewDataListViewLeftTophWidth�Height� AnchorsakLeftakTopakRightakBottom 
Checkboxes	ColumnsCaptionDataTagWidth�  CaptionPlatsWidth�  ColumnClickHideSelection
Items.Data
�   �         ��������        General configurationX   ��������        Stored sessionsX   ��������        Cached host keysX   ��������        Configuration INI fileX   ��������        Random seed fileX   ��������        Temporary foldersXReadOnly		RowSelect	ParentShowHintShowHint	TabOrder 	ViewStylevsReport	OnInfoTipDataListViewInfoTipOnKeyUpDataListViewKeyUpOnMouseDownDataListViewMouseDown  TButtonCheckAllButtonLeftTop
WidthYHeightAnchorsakLeftakBottom CaptionMarkera &allaTabOrderOnClickCheckAllButtonClick  TButton
HelpButtonLeft�TopWidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrderOnClickHelpButtonClick      TPF0TConsoleDialogConsoleDialogLeft]Top� Width7Height�HelpType	htKeywordHelpKeyword
ui_consoleBorderIconsbiSystemMenu
biMaximizebiHelp CaptionKonsolColor	clBtnFaceConstraints.MinHeight� Constraints.MinWidth|
ParentFont	OldCreateOrder	OnShowFormShow
DesignSize/� PixelsPerInch`
TextHeight TBevelBevel1Left Top Width/HeightNAlignalTopShapebsBottomLine  TLabelLabel1LeftTopWidthMHeightCaptionAnge &kommando:FocusControlCommandEdit  TLabelLabel2LeftTop8WidthPHeightCaptionAktuell katalog:  TLabelLabel4LeftTop"Width�HeightAnchorsakLeftakTopakRight AutoSizeCaptionKVarning: K�r inga kommandon som kr�ver anv�ndardata eller data�verf�ringar.  
TPathLabelDirectoryLabelLeftxTop8WidthQHeightIndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TMemo
OutputMemoLeft TopNWidth/Height?TabStopAlignalClientColor	clBtnFace	PopupMenu	PopupMenuReadOnly	
ScrollBarsssBothTabOrderWantReturnsOnContextPopupOutputMemoContextPopup  TButton	CancelBtnLeft�TopWidthKHeightAnchorsakTopakRight Cancel	CaptionSt�ngModalResultTabOrder  THistoryComboBoxCommandEditLeftxTop	Width� HeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeight	MaxLength� TabOrder OnChangeCommandEditChange  TButtonExecuteButtonLeft�TopWidthKHeightAnchorsakTopakRight CaptionK&�rDefault	TabOrderOnClickExecuteButtonClick  TButton
HelpButtonLeft�Top*WidthKHeightAnchorsakTopakRight Caption&Hj�lpTabOrderOnClickHelpButtonClick  
TImageListImagesLeft�Top� Bitmap
&  IL     �������������BM6       6   (   @                                                                                                                                                                                                                                                                                                                                                                                                                                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                                 �   �   �   �   �   �   �   �   �               �           �           �           �               ���                         �                           ���                                                                                                 �   ��� ��� ��� ��� ��� ��� ��� �       �           �           �           �           �           ���                     �   �   �                       ���                                                                                                 �   ���                     ��� �           �                                               �       ���                 �   �   �   �   �                   ���                                                                                                 �   ��� ��� ��� ��� ��� ��� ��� �               �                                   �               ���                         �                           ���                                                                             ��� ��� ��� ��� ��� �   ���                     ��� �       �                                               �           ���         �               �               �           ���                                                                             ���                 �   ��� ��� ��� ��� ��� ��� ��� �           �                                               �       ���     �   �                               �   �       ���                                                                             ��� ��� ��� ��� ��� �   ���         ��� �   �   �   �               �                                   �               ��� �   �   �   �   �               �   �   �   �   �   ���                                                                             ���                 �   ��� ��� ��� ��� �   ��� �           �                                               �           ���     �   �                               �   �       ���                                                                             ��� ��� ��� ��� ��� �   ��� ��� ��� ��� �   �                   �                                               �       ���         �               �               �           ���                                                                             ���         ���     �   �   �   �   �   �                           �                                   �               ���                         �                           ���                                                                             ��� ��� ��� ���     ���                                     �           �                                   �           ���                 �   �   �   �   �                   ���                                                                             ��� ��� ��� ���                                                 �           �           �           �           �       ���                     �   �   �                       ���                                                                                                                                                 �           �           �           �               ���                         �                           ���                                                                                                                                                                                                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                     BM>       >   (   @            �                       ��� ������  ����   � �~�  � ��|}  � ��x=  � �~�  � ��n�  � ٝO�  � ��  ��O�  �۝n�  ��7~�  ���x=  ���m|}  ���~�  ����                           
TPopupMenu	PopupMenuImagesImagesLeft�Top�  	TMenuItemCopyItemActionEditCopy  	TMenuItemSelectAllItemActionEditSelectAll  	TMenuItemN1Caption-  	TMenuItemAdjustWindowItemActionAdjustWindow   TActionList
ActionListImagesImages	OnExecuteActionListExecuteOnUpdateActionListUpdateLeft�Top�  	TEditCopyEditCopyCaptionK&opiera
ImageIndex ShortCutC@  TEditSelectAllEditSelectAllCaption&Markera allt
ImageIndexShortCutA@  TActionAdjustWindowCaptionAnpassa &F�nster
ImageIndexShortCutJ@     TPF0TCopyDialog
CopyDialogLeftkTop� HelpType	htKeywordHelpKeywordui_copyBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption
CopyDialogClientHeight� ClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameMS Sans Serif
Font.Style OldCreateOrderPositionpoMainFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize��  PixelsPerInch`
TextHeight TLabelDirectoryLabelLeftTopWidth� HeightCaption)Copy 2 selected files to remote directory  THistoryComboBoxLocalDirectoryEditLeftTopWidth�HeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeightTabOrder TextLocalDirectoryEditOnChangeControlChange  THistoryComboBoxRemoteDirectoryEditLeftTopWidth�HeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeight	MaxLength�TabOrderTextRemoteDirectoryEditOnChangeControlChange  TButton
CopyButtonLeftTop� WidthKHeightAnchorsakRightakBottom CaptionKopieraDefault	ModalResultTabOrder	  TButtonCancelButtonLeftWTop� WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder
  TButtonLocalDirectoryBrowseButtonLeft�TopWidthKHeightCaption&Bl�ddra...TabOrderOnClickLocalDirectoryBrowseButtonClick  	TCheckBoxQueueCheck2LeftTop� Width-HeightCaption1Transfer on background (add to transfer &queue) XTabOrderOnClickControlChange  	TCheckBoxQueueIndividuallyCheckLeft8Top� Width� HeightCaption'&L�gg till varje fil individuellt i k�nTabOrderOnClickControlChange  TButton
HelpButtonLeft�Top� WidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrderOnClickHelpButtonClick  	TCheckBoxNewerOnlyCheckLeftToppWidth-HeightCaptionBara &nya och �ndrade fil(er)TabOrder  	TCheckBoxNeverShowAgainCheckLeft8ToppWidth� HeightCaption#&Visa inte den h�r dialogrutan igenTabOrderOnClickControlChange  TButtonTransferSettingsButtonLeftTop� Width� HeightAnchorsakLeftakBottom Caption�verf�rin&gsinst�llningar...TabOrderOnClickTransferSettingsButtonClick  	TGroupBoxCopyParamGroupLeftTop5Width�Height2Caption�verf�ringsinst�llningarTabOrderOnContextPopupCopyParamGroupContextPopup
OnDblClickCopyParamGroupDblClick
DesignSize�2  TLabelCopyParamLabelLeftTopWidth�HeightAnchorsakLeftakTopakRightakBottom AutoSizeCaptionCopyParamLabelWordWrap	
OnDblClickCopyParamGroupDblClick      TPF0TCopyParamCustomDialogCopyParamCustomDialogLeftvTop� HelpType	htKeywordHelpKeywordui_transfer_customBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption�verf�ringsinst�llningarClientHeight�ClientWidthyColor	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameMS Sans Serif
Font.Style OldCreateOrderPositionpoMainFormCenterOnCloseQueryFormCloseQuery
DesignSizey� PixelsPerInch`
TextHeight TButtonOkButtonLeft}TopfWidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� TopfWidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  �TCopyParamsFrameCopyParamsFrameLeft Top WidthyHeightcHelpType	htKeywordTabOrder   TButton
HelpButtonLeft%TopfWidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrderOnClickHelpButtonClick     TPF0TCopyParamPresetDialogCopyParamPresetDialogLeftTopzHelpType	htKeywordHelpKeywordui_transfer_presetBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionCopyParamPresetDialogClientHeight�ClientWidthxColor	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameMS Sans Serif
Font.Style OldCreateOrderPositionpoMainFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSizex� PixelsPerInch`
TextHeight TLabelLabel1LeftTopWidthWHeightCaptionF�rinst�llnings&beskrivningFocusControlDescriptionEdit  TButtonOkButtonLeft|Top�WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft�Top�WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TEditDescriptionEditLeftTopWidthnHeight	MaxLength� TabOrder OnChangeControlChange  �TCopyParamsFrameCopyParamsFrameLeftTop3WidthyHeightcHelpType	htKeywordTabOrder  	TGroupBox	RuleGroupLeft�Top[Width� Height2AnchorsakLeftakTopakRight CaptionRegler f�r automatiskt valTabOrder
DesignSize� 2  TLabelLabel2Left
TopWidthOHeightCaptionMask v�rdna&mnFocusControlHostNameEdit  TLabelLabel3Left
TopDWidthOHeightCaptionMask an&v�ndarnamnFocusControlUserNameEdit  TLabelLabel4Left
ToptWidthoHeightCaptionMask &fj�rrkatalogFocusControlRemoteDirectoryEdit  TLabelLabel5Left
Top� WidthdHeightCaptionMask &lokal katalogFocusControlLocalDirectoryEdit  TEditHostNameEditLeft
Top$Width� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder OnChangeControlChangeOnExitMaskEditExit  TEditUserNameEditLeft
TopTWidth� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrderOnChangeControlChangeOnExitMaskEditExit  TEditRemoteDirectoryEditLeft
Top� Width� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrderOnChangeControlChangeOnExitMaskEditExit  TEditLocalDirectoryEditLeft
Top� Width� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrderOnChangeControlChangeOnExitMaskEditExit  TButtonCurrentRuleButtonLeft
Top� WidthKHeightCaptionAktuellTabOrderOnClickCurrentRuleButtonClick  TStaticTextRuleMaskHintTextLeftTop� WidthaHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaptionMasktipsTabOrderTabStop	   	TCheckBoxHasRuleCheckLeft�TopBWidth� HeightAnchorsakLeftakTopakRight Caption%V�lj automatiskt f�rinst�llningen n�rTabOrderOnClickControlChange  TButton
HelpButtonLeft$Top�WidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrderOnClickHelpButtonClick     TPF0TCopyParamsFrameCopyParamsFrameLeft Top WidthyHeightcHelpType	htKeywordTabOrder  	TGroupBoxCommonPropertiesGroupLeft� Top� Width� Height_Caption
EgenskaperTabOrder
DesignSize� _  TLabelSpeedLabel2LeftTopDWidthEHeightCaption&Hastighet (KiB/s)FocusControl
SpeedCombo  	TCheckBoxPreserveTimeCheckLeftTopWidth� HeightAnchorsakLeftakTopakRight CaptionBeh�ll tidsst�&mpelParentShowHintShowHint	TabOrder OnClickControlChange  	TCheckBoxCommonCalculateSizeCheckLeftTop,Width� HeightAnchorsakLeftakTopakRight CaptionB&er�kna total storlekParentShowHintShowHint	TabOrderOnClickControlChange  THistoryComboBox
SpeedComboLeftYTop@WidthPHeightAutoComplete
ItemHeightTabOrderText
SpeedComboOnExitSpeedComboExitItems.Strings	Unlimited10245122561286432168    	TGroupBoxLocalPropertiesGroupLeft� Top� Width� Height+Caption
EgenskaperTabOrder
DesignSize� +  	TCheckBoxPreserveReadOnlyCheckLeftTopWidth� HeightAnchorsakLeftakTopakRight CaptionBeh�ll skrivsky&ddParentShowHintShowHint	TabOrder    	TGroupBoxRemotePropertiesGroupLeftTop� Width� Height� Caption
EgenskaperTabOrder 	TCheckBoxPreserveRightsCheckLeftTopWidth� HeightCaptionS�tt fil&r�ttigheterParentShowHintShowHint	TabOrder OnClickControlChange  
TComboEdit
RightsEditLeftTop'WidthmHeight
ButtonHintKonfigurera filr�ttigheterClickKey@ParentShowHintShowHint	TabOrderText
RightsEditOnButtonClickRightsEditButtonClickOnExitRightsEditExitOnContextPopupRightsEditContextPopup  	TCheckBoxIgnorePermErrorsCheckLeftTopCWidth� HeightCaptionIgn&orera filr�ttighetsfelParentShowHintShowHint	TabOrderOnClickControlChange  	TCheckBoxClearArchiveCheckLeftTop^Width� HeightCaptionRensa 'Arki&v' attributTabOrder   	TGroupBoxChangeCaseGroupLeft� TopWidth{Height� CaptionF�r�ndra filnamnTabOrder
DesignSize{�   TRadioButtonCCLowerCaseShortButtonLeftTop^WidthnHeightAnchorsakLeftakTopakRight CaptionGemener &8.3TabOrder  TRadioButtonCCNoChangeButtonLeftTopWidthnHeightAnchorsakLeftakTopakRight CaptionI&ngen f�r�ndringTabOrder   TRadioButtonCCUpperCaseButtonLeftTop,WidthnHeightAnchorsakLeftakTopakRight Caption	&VersalerTabOrder  TRadioButtonCCLowerCaseButtonLeftTopEWidthnHeightAnchorsakLeftakTopakRight Caption&GemenerTabOrder  	TCheckBoxReplaceInvalidCharsCheckLeftTopxWidthiHeightCaptionErs�tt '\:*?' ...TabOrderOnClickControlChange   	TGroupBoxTransferModeGroupLeftTopWidth� Height� Caption�verf�ringsl�geTabOrder 
DesignSize� �   TLabelAsciiFileMaskLabelLeft
TopcWidth� HeightAnchorsakLeftakTopakRight Caption"�verf�r f�ljande &filer i textl�geFocusControlAsciiFileMaskCombo  TRadioButtonTMTextButtonLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption&Text (text, html, skript, ...)TabOrder OnClickControlChange  TRadioButtonTMBinaryButtonLeftTop0Width� HeightAnchorsakLeftakTopakRight Caption&Bin�rt (arkiv, doc, ...)TabOrderOnClickControlChange  TRadioButtonTMAutomaticButtonLeftTopJWidth� HeightAnchorsakLeftakTopakRight Caption&AutomatisktTabOrderOnClickControlChange  THistoryComboBoxAsciiFileMaskComboLeft	TopsWidth� HeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeight	MaxLength�TabOrderTextAsciiFileMaskComboOnExitValidateMaskComboExit   	TGroupBox
OtherGroupLeftTop,WidthjHeight.Caption�vrigtTabOrder
DesignSizej.  TLabelExclusionFileMaskLabelLeftZTopWidthHeightCaptionmas&k:FocusControlExcludeFileMaskCombo  THistoryComboBoxExcludeFileMaskComboLeft� TopWidth� HeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeight	MaxLength�TabOrderTextExcludeFileMaskComboOnExitValidateMaskComboExit  	TComboBoxNegativeExcludeComboLeft
TopWidthLHeightStylecsDropDownList
ItemHeightTabOrder Items.Strings	Exkludera	Inkludera    TStaticTextExcludeFileMaskHintTextLeft/TopRWidth6Height	AlignmenttaCenterCaptionMasktipsTabOrderTabStop	      TPF0TCreateDirectoryDialogCreateDirectoryDialogLeft�Top� HelpType	htKeywordHelpKeywordui_create_directoryBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption
Skapa mappClientHeight� ClientWidthQColor	clBtnFace
ParentFont	OldCreateOrder	PositionpoMainFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSizeQ�  PixelsPerInch`
TextHeight TLabel	EditLabelLeftTopWidthSHeightCaptionNytt &mappnamn:  TEditDirectoryEditLeftTopWidthAHeightAnchorsakLeftakTopakRight 	MaxLength�TabOrder TextDirectoryEditOnChangeDirectoryEditChange  TPanel	MorePanelLeft Top2WidthQHeight� AnchorsakLeftakTopakRightakBottom 
BevelOuterbvNoneTabOrder
DesignSizeQ�   	TGroupBoxAttributesGroupLeftTopWidthBHeight� AnchorsakLeftakTopakRightakBottom Caption
EgenskaperTabOrder  �TRightsExtFrameRightsFrameLeftTop$Width� HeightWTabOrder �	TCheckBoxDirectoriesXCheckVisible   	TCheckBoxSetRightsCheckLeftTopWidth� HeightCaptionS�tt fil&r�ttigheterParentShowHintShowHint	TabOrder OnClickControlChange  	TCheckBoxSaveSettingsCheckLeftTop� Width-HeightCaption&Anv�nd &samma inst�llningar n�sta g�ngTabOrder    TButtonOKBtnLeft[Top� WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeft� Top� WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeft� Top� WidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrderOnClickHelpButtonClick    TPF0TCustomCommandDialogCustomCommandDialogLeft�Top� HelpType	htKeywordHelpKeywordui_customcommandBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionCustomCommandDialogClientHeightClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameMS Sans Serif
Font.Style OldCreateOrderPositionpoMainFormCenterOnCloseQueryFormCloseQuery
DesignSize� PixelsPerInch`
TextHeight 	TGroupBoxGroupLeftTopWidth|Height� AnchorsakLeftakTopakRightakBottom TabOrder 
DesignSize|�   TLabelDescriptionLabelLeftTopWidth8HeightAnchorsakLeftakTopakRight Caption&BeskrivningFocusControlDescriptionEdit  TLabelLabel1LeftTop@WidthWHeightAnchorsakLeftakTopakRight Caption&Eget kommando:FocusControlCommandEdit  TLabelShortCutLabelLeftTop� WidthYHeightCaptionKor&tkommando:FocusControlShortCutCombo  TEditDescriptionEditLeftTop WidthfHeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder OnChangeControlChange  THistoryComboBoxCommandEditLeftTopPWidthfHeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeight	MaxLength� TabOrderOnChangeControlChange	OnGetDataCommandEditGetData	OnSetDataCommandEditSetData  	TCheckBoxApplyToDirectoriesCheckLeftTop� Width� HeightCaption&Anv�nd p� katalogerTabOrderOnClickControlChange  	TCheckBoxRecursiveCheckLeft� Top� Width� HeightCaptionK�r &rekursivtTabOrderOnClickControlChange  TRadioButtonLocalCommandButtonLeft� TopzWidth� HeightCaption&Lokalt kommandoTabOrderOnClickControlChange  TRadioButtonRemoteCommandButtonLeftTopzWidth� HeightCaption&Fj�rrkommandoTabOrderOnClickControlChange  	TCheckBoxShowResultsCheckLeftTop� Width� HeightCaption &Visa resultat i terminalf�nsterTabOrderOnClickControlChange  	TCheckBoxCopyResultsCheckLeft� Top� Width� HeightCaption&Kopiera resultat till urklippTabOrderOnClickControlChange  TStaticTextHintTextLeft"TopgWidthOHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption&m�nsterTabOrderTabStop	  	TComboBoxShortCutComboLeft� Top� Width� Height
ItemHeightTabOrder	   TButtonOkButtonLeft� Top� WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top� WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeft8Top� WidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrderOnClickHelpButtonClick   TPF0TCustomDialogCustomDialogLeft�Top� BorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSave session asXClientHeight)ClientWidthFColor	clBtnFace
ParentFont	OldCreateOrder	PositionpoMainFormCenter
DesignSizeF) PixelsPerInch`
TextHeight TButtonOKButtonLeftETop	WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top	WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder   TButton
HelpButtonLeft� Top	WidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrderOnClickHelpButtonClick   TPF0TCustomScpExplorerFormCustomScpExplorerFormLeft� Top� Width|Height�CaptionCustomScpExplorerFormColor	clBtnFace
ParentFont	
KeyPreview	OldCreateOrderPositionpoDefaultPosOnly
OnActivateFormActivateOnCloseQueryFormCloseQueryOnConstrainedResizeFormConstrainedResizeOnShowFormShowPixelsPerInch`
TextHeight 	TSplitterQueueSplitterLeft Top!WidthlHeightCursorcrVSplitHintKDra f�r att �ndra storlek p� k�listan. Dubbelklicka f�r att g�mma k�listan.AlignalBottomAutoSnapMinSizeFResizeStylersUpdateOnCanResizeQueueSplitterCanResize  TTBXDockTopDockLeft Top WidthlHeight	FixAlign	  TPanelRemotePanelLeft Top	WidthlHeightAlignalClient
BevelOuterbvNoneTabOrder  	TSplitterRemotePanelSplitterLeft� Top WidthHeightCursorcrHSplitAutoSnapMinSizeFResizeStylersUpdate  TTBXStatusBarRemoteStatusBarLeft TopWidthlHeightPanels ParentShowHintShowHint	UseSystemFontOnClickRemoteStatusBarClick  TUnixDirViewRemoteDirViewLeft� Top Width�HeightAlignalClientFullDrag	HideSelection	PopupMenu&NonVisualDataModule.RemoteDirViewPopupTabOrder	ViewStylevsReportOnColumnRightClickDirViewColumnRightClick	OnEditingDirViewEditingOnEnterRemoteDirViewEnter
NortonLikenlOffUnixColProperties.ExtWidthUnixColProperties.TypeVisibleOnDDDragFileNameRemoteFileControlDDDragFileNameOnGetSelectFilterRemoteDirViewGetSelectFilterOnLoadedDirViewLoaded
OnExecFileDirViewExecFileOnMatchMaskDirViewMatchMaskOnGetOverlayRemoteDirViewGetOverlayOnDDDragEnterFileControlDDDragEnterOnDDDragLeaveFileControlDDDragLeaveOnDDQueryContinueDrag$RemoteFileControlDDQueryContinueDragOnDDGiveFeedbackRemoteFileControlDDGiveFeedbackOnDDChooseEffectRemoteFileContolDDChooseEffectOnDDDragDetectRemoteFileControlDDDragDetectOnDDEndRemoteFileControlDDEndOnDDCreateDragFileList%RemoteFileControlDDCreateDragFileListOnDDFileOperation RemoteFileControlDDFileOperationOnDDCreateDataObject#RemoteFileControlDDCreateDataObjectOnContextPopupRemoteDirViewContextPopupOnHistoryChangeDirViewHistoryChangeOnDisplayPropertiesRemoteDirViewDisplayProperties  TUnixDriveViewRemoteDriveViewLeft Top Width� HeightDirViewRemoteDirViewOnDDDragFileNameRemoteFileControlDDDragFileNameOnDDEndRemoteFileControlDDEndUseSystemContextMenuOnDDDragEnterFileControlDDDragEnterOnDDDragLeaveFileControlDDDragLeaveOnDDQueryContinueDrag$RemoteFileControlDDQueryContinueDragOnDDChooseEffectRemoteFileContolDDChooseEffectOnDDGiveFeedbackRemoteFileControlDDGiveFeedbackOnDDDragDetectRemoteFileControlDDDragDetectOnDDFileOperation RemoteFileControlDDFileOperationOnDDCreateDragFileList%RemoteFileControlDDCreateDragFileListOnDDCreateDataObject#RemoteFileControlDDCreateDataObjectAlignalLeftIndentParentColorReadOnly	TabOrderOnEnterRemoteDriveViewEnter   TPanel
QueuePanelLeft Top$WidthlHeight� AlignalBottom
BevelOuterbvNoneTabOrder 	TListView
QueueView2Left TopWidthlHeightrAlignalClientColumnsCaption	OperationWidthF CaptionK�llaWidth�  CaptionM�lWidth�  	AlignmenttaRightJustifyCaption�verf�rtWidthP 	AlignmenttaRightJustifyCaptionTid/HastighetWidthP 	AlignmenttaCenterCaption
UtvecklingWidthP  ColumnClickDragModedmAutomaticReadOnly		RowSelect		PopupMenuNonVisualDataModule.QueuePopupSmallImagesGlyphsModule.QueueImagesStateImagesGlyphsModule.QueueImagesTabOrder 	ViewStylevsReportOnContextPopupQueueView2ContextPopup
OnDeletionQueueView2DeletionOnEnterQueueView2Enter
OnDragDropQueueView2DragDrop
OnDragOverQueueView2DragOverOnSelectItemQueueView2SelectItemOnStartDragQueueView2StartDrag  TTBXDock	QueueDockTagLeft Top WidthlHeight	AllowDrag TTBXToolbarQueueToolbarLeft Top CaptionQueueToolbarImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder  TTBXItem
TBXItem201Action(NonVisualDataModule.QueueItemQueryAction  TTBXItem
TBXItem202Action(NonVisualDataModule.QueueItemErrorAction  TTBXItem
TBXItem203Action)NonVisualDataModule.QueueItemPromptAction  TTBXItem
TBXItem204Action*NonVisualDataModule.QueueItemExecuteAction  TTBXItem
TBXItem195Action(NonVisualDataModule.QueueItemPauseAction  TTBXItem
TBXItem194Action)NonVisualDataModule.QueueItemResumeAction  TTBXItem
TBXItem205Action)NonVisualDataModule.QueueItemDeleteAction  TTBXSeparatorItemTBXSeparatorItem201  TTBXItem
TBXItem206Action%NonVisualDataModule.QueueItemUpAction  TTBXItem
TBXItem207Action'NonVisualDataModule.QueueItemDownAction  TTBXSeparatorItemTBXSeparatorItem202  TTBXSubmenuItemTBXSubmenuItem27Action-NonVisualDataModule.QueueCycleOnceEmptyActionDropdownCombo	 TTBXItem
TBXItem211Action,NonVisualDataModule.QueueIdleOnceEmptyAction	RadioItem	  TTBXItem
TBXItem225Action2NonVisualDataModule.QueueDisconnectOnceEmptyAction	RadioItem	  TTBXItem
TBXItem226Action0NonVisualDataModule.QueueShutDownOnceEmptyAction	RadioItem	   TTBXItem
TBXItem208Action*NonVisualDataModule.QueuePreferencesAction       TPF0TEditorForm
EditorFormLeft;Top� WidthqHeight�HelpType	htKeywordHelpKeyword	ui_editorBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp Caption
EditorFormColor	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameMS Sans Serif
Font.Style 	Icon.Data
>           (     (                �                         �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                 x�����  �����  x����  ��� �  ���    ����  ���x0  �����  ����  ����;0 ��� 8� ���� ���p� wwwwp  ��                                          !   s  
KeyPreview	OldCreateOrderPositionpoDefaultPosOnly
OnActivateFormActivateOnClose	FormCloseOnCloseQueryFormCloseQueryOnShowFormShowPixelsPerInch`
TextHeight TTBXDockTopDockLeft Top WidthiHeight	AllowDrag TTBXToolbarToolBarLeft Top CaptionToolBarImagesEditorImagesParentShowHintShowHint	TabOrder  TTBXItemTBXItem1ActionCloseAction  TTBXItemTBXItem2Action
SaveAction  TTBXItem	TBXItem16ActionReloadAction  TTBXSeparatorItemTBXSeparatorItem1  TTBXItemTBXItem3ActionEditCopy  TTBXItemTBXItem4ActionEditCut  TTBXItemTBXItem5Action	EditPaste  TTBXItemTBXItem6Action
EditDelete  TTBXItemTBXItem7ActionEditSelectAll  TTBXSeparatorItemTBXSeparatorItem2  TTBXItemTBXItem8ActionEditUndo  TTBXItem	TBXItem17ActionEditRedo  TTBXSeparatorItemTBXSeparatorItem3  TTBXItemTBXItem9Action
FindAction  TTBXItem	TBXItem10ActionReplaceAction  TTBXItem	TBXItem11ActionFindNextAction  TTBXItem	TBXItem12ActionGoToLineAction  TTBXSeparatorItemTBXSeparatorItem4  TTBXItem	TBXItem13ActionPreferencesAction  TTBXSeparatorItemTBXSeparatorItem5  TTBXItem	TBXItem14Action
HelpAction    TTBXStatusBar	StatusBarLeft TopkWidthiPanelsCaptionLine: 2000/20000Size� Tag  Caption
Column: 20ViewPriorityPSize� Tag  CaptionCharacter: 132 (0x56)ViewPriorityZSize� Tag  ViewPriorityFStretchPrioritydTag   UseSystemFont  TActionListEditorActionsImagesEditorImages	OnExecuteEditorActionsExecuteOnUpdateEditorActionsUpdateLeft�Top8 TAction
SaveActionCaption&SparaHintSpara|Spara fil
ImageIndex ShortCutS@SecondaryShortCuts.StringsF2   TEditCutEditCutCaption
K&lipp u&tHint?Klipp ut|Klipper ut vald markering och flyttar det till urklipp
ImageIndexShortCutX@  	TEditCopyEditCopyCaption&KopieraHint,Kopiera|Kopierar vald markering till urklipp
ImageIndexShortCutC@  
TEditPaste	EditPasteCaptionKl&istra inHint.Klistra in|Klistrar in inneh�llet fr�n urklipp
ImageIndexShortCutV@SecondaryShortCuts.Strings	Shift+InsCtrl+Shift+Ins   TEditSelectAllEditSelectAllCaptionM&arkera alltHint%Markera allt|Markerar hela dokumentet
ImageIndexShortCutA@  	TEditUndoEditUndoCaption&�ngraHint"�ngra|�ngrar den senaste �ndringen
ImageIndexShortCutZ@  TActionEditRedoCaption&G�r omHint#G�r om|G�r om den senaste �ndringen
ImageIndexShortCutY@  TEditDelete
EditDeleteCaption&RaderaHintRadera|Raderar vald markering
ImageIndex  TActionPreferencesActionCaption&Inst�llningar...Hint7Inst�llningar|Visa/�ndra textredigerarens inst�llningar
ImageIndex  TActionCloseActionCaptionS&t�ngHint9St�ng|Spara filen om n�dv�ndigt och st�ng textredigeraren
ImageIndexShortCut  TAction
FindActionCaption&S�k...HintS�k|S�k den valda texten
ImageIndex	ShortCutF@SecondaryShortCuts.StringsF7   TActionReplaceActionCaption
&Ers�tt...Hint0Ers�tt|Ers�tt den valda texten med en annan text
ImageIndex
ShortCutH@SecondaryShortCuts.StringsCtrl+F7   TActionFindNextActionCaption
S�k &n�staHint6S�k n�sta|S�k efter n�sta uppkomst av den valda texten
ImageIndexShortCutrSecondaryShortCuts.StringsShift+F7   TActionGoToLineActionCaption&G� till radnummer...Hint-G� till radnummer|G� till det valda radnumret
ImageIndexShortCutG@SecondaryShortCuts.StringsAlt+F8   TAction
HelpActionCaption&Hj�lpHintHj�lp editor
ImageIndex  TActionReloadActionCaption	La&dda omHintLadda om|Laddar om fil
ImageIndexShortCutR@   
TImageListEditorImagesLeftTop8Bitmap
&S  IL     �������������BM6       6   (   @   P           P                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                               �                       �   �   �   �   �                                                                                                                                                                                                                   �                               �   �   �   �                                                                                                                                                                                                                   �                                   �   �   �                                                                                                                                                                                                                   �                               �       �   �                                                                                                                                                                                                                       �                   �   �               �                                                                                                                                                                                                                           �   �   �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               f f                                                                                                                                                                                 ���                                                                 f f f f � � � �                                                                                                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 f f f f � � �f� ��� ��� � �                                                                                             ��� ��� ��� ��� ��� ���  �1 ��� ��� ��� ��� ���                             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���         f f f f � � �f� ��� ��� ��� ��� ��� � �                                                             �   �   �                   ��� ��� ��� ��� ���  �1  �1 ��� ��� ��� ��� ���             �               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���     � � � � �f� ��� ��� ��� ��� � � ��� ��� ��� � �                                                         �   �   �                   ��� ��� ��� ���  �1  �1  �1  �1  �1 ��� ��� ���             �   �           ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���     � � ��� ��� ��� ��� � � � � � �     ��� ��� ��� � �                                                                                 ��� ��� ��� ��� ���  �1  �1 ��� c�  cc  ��� ���             �   �   �       ���  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��     � � ��� ��� � � � � � � � � � � � �     fff ��� ��� � �                                                 �   �   �                   ��� ��� ��� ��� ��� ���  �1 ��� ��� cc  ��� ���             �   �   �       ���  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��     � � � � � � � � � � � � � � � � � � � �     fff ��� ��� � �                                             �   �   �                   ��� ��� ��� cc  ��� ��� ��� ��� ��� cc  ��� ���             �   �           ���  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��     � � ��� � � � � � �  �� 3�� 3f� � � � � � �     fff ��� � �                                                 �   �   �               ��� ��� ��� cc  ��� ���  �1 ��� ��� ��� ��� ���             �               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���         � � ��� � � � � � � � �  ��  �� 3�� 3f� � �     fff � � ���                                                 �   �   �           ��� ��� ��� cc  c�  ���  �1  �1 ��� ��� ��� ���                             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���             � � ��� � � � � � � � � � � 3��  �� f f � �     � � ���                             �   �   �               �   �   �       ��� ��� ��� ���  �1  �1  �1  �1  �1 ��� ��� ���                             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 � � ��� � � � �  ��  ��  �� 3�� f f � � � �                                     �   �   �               �   �   �       ��� ��� ��� ��� ��� ���  �1  �1 ��� ��� ��� ���                             ��� ��� ��� ��� ��� ��� ��� ���                                 � � ��� � � � � 3f� 3f� f f � � � � f f                                     �   �   �               �   �   �       ��� ��� ��� ��� ��� ���  �1 ��� ���                                         ��� ��� ��� ��� ��� ��� ��� ���     ���                             � � ��� � � � � � � � � f f                                                 �   �   �   �   �   �   �           ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                 ��� ��� ��� ��� ��� ��� ��� ���                                         � � ��� � � f f                                                             �   �   �   �   �               ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                     ��� ��� ��� ��� ��� ��� ��� ���                                             � �                                                                                                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                                                                                                                                                                                                                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���     ���     ���                                                                                                                                                                                                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                                                                                                                                 �   �   �   �           ��� ��� ��� ��� ��� ��� �   �   �   �       ���                                     ���                                                                                                                                                             �   �   �           ��� ��� ��� ��� �                   ���                                     ���                                                                                                                                                             �   �   �   �       ��� ��� ��� ��� �                                                                                                                                                                                                                           �   �   �   �       ��� ��� ��� ��� �                       ���                         ���                                                                                                     ���                             ���                             �   �   �   �       ��� ��  ��� ��  �                       ���             ���         ���                                     ���                             ���                                     ���             ���                                     �   �   �   �       ��  ��� ��  ��� �                       ���             ���         ���                                             ���             ���                                                                                                     �   �   �   �       ��� ��  ��� ��  �                                                                                                                                                           ���                 ���                                         �   �   �   �       ��  ��� ��  ��� �                           ���                     ���                                     ���                 ���                                         ���                 ���                                         �   �   �   �   �   �   �   �   �   �                                                                                           ���                 ���                                                                                                                                                                                                                                                                                                                         ���                                                                                                                 ���                     ���                                                 ���                                                                                                                          �   �   �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��� ��� ��� ���                                                                                                                                                                     �           �           �           �                               ���                 ���     ���                                                                                                                                                     �           �           �           �           �                               ���                 ���     ���                                                                                                                                                     �                                               �                                                           ���                                                         �                                                                                           �                                   �                       ���                                                             �   �   �   �   �                       �                                                                                   �                                               �           ��� ���                                             ��� ���             �   �   �   �                               �                                                                                   �                                               �       ���                     ��� ��� ���                                     �   �   �                                   �                                                                                       �                                   �               ���                     ��� ��� ���                                     �   �       �                               �                                                                               �                                               �           ���                     ��� ��� ���                                     �               �   �                   �                                                                                       �                                               �               ���                                                                                     �   �   �   �                                                                                               �                                   �                                                                   ���                                                                                                                                             �           �                                   �                   ���                                                                                                                                                                                             �           �           �           �           �                   ���     ���                 ���                                                                                                                                                                 �           �           �           �                                                   ���                                                                                                                                                                                                                                                 ��� ��� ��� ���                                                                                                                                                                                                                                                                                                                                                                             �   �                                                                                                                               �   �   �   �   �   �   �   �   �   �       ��� �II �NN �GG ��� ��� ��� ��� ��� ��� �44 �44 �NN �NN                     �           �           �   �                                               �   �   �   �   �   �   �   �   �                           �   ��� ��� ��� ��� ��� ��� ��� ��� �       ��v �gg �gg �NN ��� �vv ڴ� ��� ��� ��� �44 �44 �gg �NN                     �           �       �           �                                           �   ��� ��� ��� ��� ��� ��� ��� �       ���  �� ���  �� ��� �   ���                         ��� �       ��v �gg �gg �NN ϶� �RR ��� ��� ��� ��� �44 �44 �gg �NN                     �           �       �           �                                           �   ���                     ��� �        �� ���  �� ���  �� �   ��� ��� ��� ��� ��� ��� ��� ��� �       ��v �gg �gg �NN ��� �CC �ww ��� ��� ��� �44 �44 �gg �NN                         �   �   �       �           �                                           �   ��� ��� ��� ��� ��� ��� ��� �       ���  �� ���  �� ��� �   ���             ��� �   �   �   �       ��v �gg �gg �NN ��� ʗ� ʱ� ��� ��� ��� �44 �77 �gg �NN                                 �       �   �   �                           ��� ��� ��� ��� ��� �   ���                     ��� �        �� ���  �� ���  �� �   ��� ��� ��� ��� ��� �   ��� �           ��v �gg �gg �gg �gg �gg �gg �gg �gg �gg �gg �gg �gg �NN                                 �       �                                   ���                 �   ��� ��� ��� ��� ��� ��� ��� �       ���  �� ���  �� ��� �   ��� ��� ��� ��� ��� �   �               ��v �gg �gg ��� ��� ��� ��� ��� ��� ��� ��� �gg �gg �NN                                                                             ��� ��� ��� ��� ��� �   ���         ��� �   �   �   �        �� ���  �� ���  �� �   �   �   �   �   �   �                   ��v �gg ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �gg �NN                                                                             ���                 �   ��� ��� ��� ��� �   ��� �           ���  �� ���  �� ���  �� ���  �� ���  �� ���  ��                 ��v �gg ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �gg �NN                                                                             ��� ��� ��� ��� ��� �   ��� ��� ��� ��� �   �                �� ���                                 ��� ���                 ��v �gg ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �gg �NN                                                                             ���         ���     �   �   �   �   �   �                   ��� ���                                 ���  ��                 ��v �gg ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �gg �NN                                                                             ��� ��� ��� ���     ���                                      �� ���  ��      ��          ��     ���  �� ���                 ��v �gg ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �gg �NN                                                                             ��� ��� ��� ���                                                                  ��  ��                                     ��v �NN ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �NN ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                     BM>       >   (   @   P         �                      ��� ��      ��      ��      ��      ��      ��      �      ��      ��      ��      �;      ��      ��      ��      ��      ��      ������� �?���� ����� ��ǀp  sǀ0  '��  ǀ    ǀ0   �p � �� � 8�� � 8�� �8���?������������������ ���k�I  ��'�I  ��k�������������� ����� ��Ç� Ç����������������������������������������������?������/�����������������������繛 ����ٝ ���� ���?� ���۝�����7������������m�������?�������?��������������� ���� � ����   ����   ����   ����  ��?�  ���  ��?� ���� ����À�߀ ��߀����߁����������                        TTBXPopupMenuEditorPopupImagesEditorImagesLeft�Top�  TTBXItemUndo1ActionEditUndo  TTBXItem	TBXItem18ActionEditRedo  TTBXSeparatorItemN1  TTBXItemCut1ActionEditCut  TTBXItemCopy1ActionEditCopy  TTBXItemPaste1Action	EditPaste  TTBXItemDelete1Action
EditDelete  TTBXSeparatorItemN2  TTBXItem
SelectAll1ActionEditSelectAll  TTBXSeparatorItemN3  TTBXItemFind1Action
FindAction  TTBXItemReplace1ActionReplaceAction  TTBXItem	Findnext1ActionFindNextAction  TTBXItemGotolinenumber1ActionGoToLineAction  TTBXSeparatorItemTBXSeparatorItem6  TTBXItem	TBXItem15ActionPreferencesAction      TPF0TEditorPreferencesDialogEditorPreferencesDialogLeft/Top� HelpType	htKeywordHelpKeywordui_editor_preferencesBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionEditorPreferencesDialogClientHeightgClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameMS Sans Serif
Font.Style OldCreateOrderPositionpoMainFormCenterOnCloseQueryFormCloseQuery
DesignSize�g PixelsPerInch`
TextHeight 	TGroupBoxExternalEditorGroupLeftTop� Width�HeightIAnchorsakLeftakTopakRight CaptionAAlternativ extern editor (p�verkar bara redigering av fj�rrfiler)TabOrder 	TCheckBoxExternalEditorTextCheckLeftTop-WidthQHeightCaptionDTvinga fram text�verf�ringsl�ge f�r filer redigerade i extern editorTabOrder  	TCheckBoxSDIExternalEditorCheckLeftTopWidthQHeightCaption?E&xtern editor �ppnar varje fil i ett separat f�nster (process)TabOrder    	TGroupBoxEditorGroup2LeftTopWidth�Height}AnchorsakLeftakTopakRight CaptionEditorTabOrder 
DesignSize�}  TRadioButtonEditorInternalButtonLeftTopWidth� HeightCaption&Intern editorTabOrder OnClickControlChange  TRadioButtonEditorExternalButtonLeftTop-Width� HeightCaption&Extern editorTabOrderOnClickControlChange  THistoryComboBoxExternalEditorEditLeft TopEWidthHeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeightTabOrderTextExternalEditorEditOnChangeControlChangeOnExitExternalEditorEditExit  TButtonExternalEditorBrowseButtonLeft1TopCWidthKHeightCaptionB&l�ddra...TabOrderOnClickExternalEditorBrowseButtonClick  TRadioButtonEditorOpenButtonLeftTopaWidth� HeightCaption&Associerad applikationTabOrderOnClickControlChange   	TGroupBox	MaskGroupLeftTop� Width�HeightIAnchorsakLeftakTopakRight CaptionAutomatiskt val av editorTabOrder
DesignSize�I  TLabel	MaskLabelLeftTopWidth� HeightCaption+Anv�nd den h�r editorn f�r &f�ljande filer:FocusControlMaskEdit  THistoryComboBoxMaskEditLeftTop'WidthoHeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeight	MaxLength�TabOrder Text*.*OnExitMaskEditExit   TButtonOkButtonLeft� TopFWidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� TopFWidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeft?TopFWidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrderOnClickHelpButtonClick  	TCheckBoxRememberCheckLeftTop.WidthQHeightAnchorsakLeftakBottom Caption&Kom ih�g den h�r editornTabOrder      TPF0TFileFindDialogFileFindDialogLeftoTop� WidthBHeight�HelpType	htKeywordHelpKeywordui_findBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp CaptionFindXColor	clBtnFaceConstraints.MinHeight� Constraints.MinWidth^Font.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameMS Sans Serif
Font.Style 
KeyPreview	OldCreateOrderPositionpoMainFormCenterOnCloseQueryFormCloseQuery	OnKeyDownFormKeyDownOnShowFormShow
DesignSize:� PixelsPerInch`
TextHeight 	TGroupBoxFilterGroupLeftTopWidth�HeightAnchorsakLeftakTopakRight CaptionFilterTabOrder 
DesignSize�  TLabel	MaskLabelLeftTopWidth/HeightCaption	&Filmask:FocusControlMaskEdit  TLabelRemoteDirectoryLabelLeftTopGWidth0HeightCaptionS�&k i:FocusControlRemoteDirectoryEdit  THistoryComboBoxRemoteDirectoryEditLeftTopWWidth�HeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeight	MaxLength�TabOrderTextRemoteDirectoryEditOnChangeControlChange  THistoryComboBoxMaskEditLeftTop$Width�HeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeight	MaxLength�TabOrder TextMaskEditOnChangeControlChangeOnExitMaskEditExit  TStaticTextMaskHintTextLeftgTop@WidthaHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption	Mask&tipsTabOrderTabStop	   TButtonCancelButtonLeft�Top+WidthPHeightAnchorsakTopakRight Cancel	CaptionSt�ngModalResultTabOrder  TButtonStartStopButtonLeft�TopWidthPHeightAnchorsakTopakRight Caption&StartXDefault	TabOrderOnClickStartStopButtonClick  TButton
HelpButtonLeft�TopKWidthPHeightAnchorsakTopakRight Caption&Hj�lpTabOrderOnClickHelpButtonClick  TIEListViewFileViewLeftTop� Width�Height� AnchorsakLeftakTopakRightakBottom ColumnClickFullDrag	ReadOnly		RowSelect	TabOrder	ViewStylevsReport
OnDblClickFileViewDblClick
NortonLikenlOffColumnsCaptionNamnWidthP CaptionKatalogWidthx 	AlignmenttaRightJustifyCaptionStorlekWidthP Caption�ndradWidthZ  MultiSelectOnSelectItemFileViewSelectItem  
TStatusBar	StatusBarLeft Top�Width:HeightPanels ParentShowHintShowHint	SimplePanel	  TButtonFocusButtonLeft�Top� WidthPHeightAnchorsakTopakRight CaptionF&okusModalResultTabOrderOnClickFocusButtonClick  TButtonMinimizeButtonLeft�Top+WidthPHeightAnchorsakTopakRight Caption	&MinimeraTabOrderOnClickMinimizeButtonClick     TPF0TFileSystemInfoDialogFileSystemInfoDialogLeft� TopEHelpType	htKeywordHelpKeyword	ui_fsinfoBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption#Information om server och protokollClientHeightrClientWidthsColor	clBtnFace
ParentFont	OldCreateOrder	PositionpoMainFormCenterOnShowFormShow
DesignSizesr PixelsPerInch`
TextHeight TButtonCloseButtonLeft� TopPWidthKHeightAnchorsakRightakBottom Cancel	CaptionSt�ngDefault	ModalResultTabOrder  TButton
HelpButtonLeftTopPWidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrderOnClickHelpButtonClick  TPageControlPageControlLeft Top WidthsHeightD
ActivePageProtocolSheetAlignalTopAnchorsakLeftakTopakRightakBottom TabIndex TabOrder OnChangePageControlChange 	TTabSheetProtocolSheetCaption	Protokoll
DesignSizek(  	TGroupBoxHostKeyGroupLeftTop� Width_Height)AnchorsakLeftakRightakBottom Caption#Nyckelfingeravtryck till v�rdserverTabOrder
DesignSize_)  TEditHostKeyFingerprintEditLeft
TopWidthNHeightTabStopAnchorsakLeftakTopakRight BorderStylebsNoneColor	clBtnFaceReadOnly	TabOrder TextHostKeyFingerprintEdit   	TListView
ServerViewLeftTopWidth_Height� AnchorsakLeftakTopakRightakBottom ColumnsCaptionArtikelWidth�	WidthType�  CaptionV�rdeWidth�	WidthType�   ColumnClickMultiSelect	ReadOnly		RowSelect		PopupMenuListViewMenuTabOrder 	ViewStylevsReportOnContextPopupControlContextPopup  	TGroupBoxCertificateGroupLeftTop� Width_HeightHAnchorsakLeftakRightakBottom CaptionCertifikatets fingeravtryckTabOrder
DesignSize_H  TEditCertificateFingerprintEditLeft
TopWidthNHeightTabStopAnchorsakLeftakTopakRight BorderStylebsNoneColor	clBtnFaceReadOnly	TabOrder TextCertificateFingerprintEdit  TButtonCertificateViewButtonLeft
Top%WidthyHeightCaption&Fullst�ndigt certifikatTabOrderOnClickCertificateViewButtonClick    	TTabSheetCapabilitiesSheetCaptionM�jligheter
ImageIndex
DesignSizek(  	TGroupBox	InfoGroupLeftTop� Width_HeightrAnchorsakLeftakRightakBottom Caption�vrig informationTabOrder
DesignSize_r  TMemoInfoMemoLeft	TopWidthMHeightWTabStopAnchorsakLeftakTopakRight 
BevelInnerbvNone
BevelOuterbvNoneBorderStylebsNoneColor	clBtnFaceLines.StringsInfoMemo ReadOnly	
ScrollBarsssBothTabOrder WantReturnsWordWrap   	TListViewProtocolViewLeftTopWidth_Height� AnchorsakLeftakTopakRightakBottom ColumnsCaptionArtikelWidth�	WidthType�  CaptionV�rdeWidth�	WidthType�   ColumnClickMultiSelect	ReadOnly		RowSelect		PopupMenuListViewMenuTabOrder 	ViewStylevsReportOnContextPopupControlContextPopup   	TTabSheetSpaceAvailableSheetCaptionTillg�ngligt utrymme
ImageIndex
DesignSizek(  TLabelLabel1LeftTopWidthHeightCaption&S�kv�g:FocusControlSpaceAvailablePathEdit  	TListViewSpaceAvailableViewLeftTop(Width_HeightAnchorsakLeftakTopakRightakBottom ColumnsCaptionArtikelWidth�	WidthType�  CaptionV�rdeWidth�	WidthType�   ColumnClickMultiSelect	ReadOnly		RowSelect		PopupMenuListViewMenuTabOrder	ViewStylevsReportOnContextPopupControlContextPopup  TEditSpaceAvailablePathEditLeft8Top	Width� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder OnChangeControlChangeOnEnterSpaceAvailablePathEditEnterOnExitSpaceAvailablePathEditExit  TButtonSpaceAvailableButtonLeft TopWidthcHeightAnchorsakTopakRight CaptionKon&trolleraTabOrderOnClickSpaceAvailableButtonClick    TButtonClipboardButtonLeftTopPWidthyHeightAnchorsakRightakBottom Caption&Kopiera till urklippTabOrderOnClickClipboardButtonClick  
TPopupMenuListViewMenuLeft� TopH 	TMenuItemCopyCaptionK&opieraOnClick	CopyClick    TPF0TFullSynchronizeDialogFullSynchronizeDialogLeftmTop� HelpType	htKeywordHelpKeywordui_synchronizeBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSynkroniseraClientHeight�ClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameMS Sans Serif
Font.Style OldCreateOrderPositionpoMainFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize�� PixelsPerInch`
TextHeight 	TGroupBoxDirectoriesGroupLeftTopWidth�HeightwAnchorsakLeftakTopakRight Caption	KatalogerTabOrder 
DesignSize�w  TLabelLocalDirectoryLabelLeftTopWidthHHeightAnchorsakLeftakTopakRight CaptionL&okal katalog:FocusControlLocalDirectoryEdit  TLabelRemoteDirectoryLabelLeftTopDWidthSHeightAnchorsakLeftakTopakRight CaptionF&j�rrka&talog:FocusControlRemoteDirectoryEdit  THistoryComboBoxRemoteDirectoryEditLeftTopTWidth�HeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeight	MaxLength�TabOrderTextRemoteDirectoryEditOnChangeControlChange  THistoryComboBoxLocalDirectoryEditLeftTop#Width8HeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeight	MaxLength�TabOrder TextLocalDirectoryEditOnChangeControlChange  TButtonLocalDirectoryBrowseButtonLeftJTop!WidthKHeightAnchorsakTopakRight CaptionBl&�ddra...TabOrderOnClickLocalDirectoryBrowseButtonClick   TButtonOkButtonLeft� Top�WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeftTop�WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder	  	TGroupBoxOptionsGroupLeftTop� WidthHeightICaptionAlternativ f�r synkroniseringTabOrder 	TCheckBoxSynchronizeDeleteCheckLeftTopWidth~HeightCaption&Ta bort filerTabOrder OnClickControlChange  	TCheckBoxSynchronizeSelectedOnlyCheckLeft� Top,Width{HeightCaptionBara &valda filerTabOrderOnClickControlChange  	TCheckBoxSynchronizeExistingOnlyCheckLeft� TopWidth{HeightCaption&Endast existerande filerTabOrderOnClickControlChange  	TCheckBoxSynchronizePreviewChangesCheckLeftTop,Width~HeightCaptionF�&rhandsvisa �ndringarTabOrderOnClickControlChange   TButtonTransferSettingsButtonLeftTop�Width� HeightAnchorsakLeftakBottom Caption�verf&�ringsinst�llningar...TabOrderOnClickTransferSettingsButtonClick  	TGroupBoxDirectionGroupLeftTop� Width�Height1AnchorsakLeftakTopakRight CaptionRiktning/m�lkatalogTabOrder TRadioButtonSynchronizeBothButtonLeftTopWidthfHeightCaption&B�daTabOrder OnClickControlChange  TRadioButtonSynchronizeRemoteButtonLeft� TopWidthfHeightCaption&Fj�rrTabOrderOnClickControlChange  TRadioButtonSynchronizeLocalButtonLeftTopWidth� HeightCaption&LokalTabOrderOnClickControlChange   	TGroupBoxCompareCriterionsGroupLeftTop� Width� HeightICaptionJ�mf�relsekriterierTabOrder 	TCheckBoxSynchronizeByTimeCheckLeftTopWidthyHeightCaption�&ndringstidTabOrder OnClickControlChange  	TCheckBoxSynchronizeBySizeCheckLeftTop,WidthyHeightCaptionF&ilstorlekTabOrderOnClickControlChange   	TCheckBoxSaveSettingsCheckLeftTop=Width� HeightCaptionAnv�nd &samma val n�sta g�ngTabOrder  	TGroupBoxCopyParamGroupLeftTopRWidth�Height2Caption�verf�ringsinst�llningarTabOrderOnContextPopupCopyParamGroupContextPopup
OnDblClickCopyParamGroupDblClick
DesignSize�2  TLabelCopyParamLabelLeftTopWidth�HeightAnchorsakLeftakTopakRightakBottom AutoSizeCaptionCopyParamLabelWordWrap	
OnDblClickCopyParamGroupDblClick   TButton
HelpButtonLeft]Top�WidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrder
OnClickHelpButtonClick  	TGroupBox	ModeGroupLeftTop� Width�Height1AnchorsakLeftakTopakRight CaptionMetodTabOrder TRadioButtonSynchronizeFilesButtonLeftTopWidth~HeightCaptionSynkronisera &filerTabOrder OnClickControlChange  TRadioButtonMirrorFilesButtonLeft� TopWidth� HeightCaptionS&pegelfilerTabOrderOnClickControlChange  TRadioButtonSynchronizeTimestampsButtonLeftTopWidth� HeightCaptionSynkronisera tidss&t�mplarTabOrderOnClickControlChange      TPF0TGeneralSettingsFrameGeneralSettingsFrameLeft Top Width2Height� TabOrder 
DesignSize2�   	TGroupBoxInterfaceGroupLeft Top Width2Height� AnchorsakLeftakTopakRightakBottom Caption
Gr�nssnittTabOrder 
DesignSize2�   TLabelCommanderDescriptionLabel2Left� TopWidth� HeightsAnchorsakLeftakTopakRight AutoSizeCaption�- tv� paneler (v�nster f�r lokal katalog, h�ger f�r fj�rrkatalog)
- snabbkommandon som i Norton Commander (och andra liknande program som Total Commander, Midnight Commander...)
- dra && sl�pp till/fr�n b�da panelernaWordWrap	OnClickCommanderClick  TLabelExplorerDescriptionLabelLeft� Top� Width� Height>AnchorsakLeftakTopakRight AutoSizeCaptionI- endast fj�rrkatalog
- snabbkommandon som i Utforskaren
- dra && sl�ppWordWrap	OnClickExplorerClick  TImageCommanderInterfacePictureLeft7Top)Width Height AutoSize	Picture.Data
B  TBitmap6  BM6      6   (                    �  �                                                                                                          ���������������������������������������������������������������������������������������������   �����������������������������������������������������������������������������������������Ƅ��   ������      ��ƀ�����������������      ��ƀ�����������������      ��ƀ�������������������Ƅ��   �����Ƅ����������������������������������������������������������������������������������Ƅ��   �����������������������������������������������������������������������������������������Ƅ��   ��������� �  � ��������������������������������������������������������������������������Ƅ��   �������������  ���      ������������      �����������������������������������������������Ƅ��   �����������������������������������������������������������������������������������������Ƅ��   ����������  � ���������������������������������������������������������������������������Ƅ��   ������������� ����            ������      �����������������������������������������������Ƅ��   �����������������������������������������������������������������������������������������Ƅ��   ��������� � �  ������������������������������������� ��  ��������������������������������Ƅ��   �������������  ���         ���������      ������������� ����         ���������      �����Ƅ��   �����������������������������������������������������������������������������������������Ƅ��   ����������    ��������������������������������������  �� ��������������������������������Ƅ��   �������������  ���               ���      �������������  ���               ���      �����Ƅ��   �����������������������������������������������������������������������������������������Ƅ��   ��������� ���  ������������������������������������ ���  ��������������������������������Ƅ��   ������������ �����            ������      ������������ �����            ������      �����Ƅ��   �����������������������������������������������������������������������������������������Ƅ��   �����Ƅ����������������������������������������������������������������������������������Ƅ��   �����Ƅ����� �� � ��� ���  ���@���� @@ ���  �� ���ƀ� � ����@��� �  ���������������������Ƅ��   �����Ƅ�� �����  �����  ��ƀ ������ƀ ��� ��ƀ�  �������� @���� � ����� �����������������Ƅ��   �����Ƅ����������������������������������������������������������������������������������Ƅ��   �����������������������������������������������������������������������������������������Ƅ��   �����Ƅ  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �                             ���   �����Ƅ  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ������   ������   ������   ���   �����Ƅ  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ������   ������   ������   ���   �����Ƅ  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ���   �����������������������������������������������������������������������������������������Ƅ��   ���������������������������������������������������������������������������������������������   OnClickCommanderClick  TImageExplorerInterfacePictureLeft7Top� Width Height AutoSize	Picture.Data
B  TBitmap6  BM6      6   (                    �  �          ����������                                                                                 ����������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������Ƅ��   ������������������������������������������������������������������������������������Ƅ��   ����������������������      �� ������������@@ � @@@ ��������������������������������Ƅ��   ������������������������ �� �� ������������@��� @@@ ��������������������������������Ƅ��   �����������������������   �    ������������@��@��@����������������������������������Ƅ��                  ��������������������������������������������������������������������������Ƅ��   �����������������������������������������������������������������������������������������Ƅ��   ��������������Ƅ�������������������������������������������������������������������������Ƅ��   ��������������������������� � � �� ������������� � � �� @������������� ���    �����������Ƅ��   ������������   ������������ �    � ������������� � � �� @������������� ���    �����������Ƅ��   �������������� ������������ �� �    �������������� �� � @������������� ��� �� �����������Ƅ��   �������������  ��������������������������������������������������������������������������Ƅ��   ��������������������Ƅ�������������������������������������������������������������������Ƅ��   ��������������������Ƅ����� �� � ��� ���  ���@���� @@ � ����@��� �  ���������������������Ƅ��   ��������������������Ƅ�� �����  �����  ��ƀ ������ƀ ���� @���� � ����� �����������������Ƅ��   ������������ � �����Ƅ�������������������������������������������������������������������Ƅ��   ������������ � ��������������������������������������������������������������������������Ƅ��   ������������ �������Ƅ  �  �  �  �  �  �  �  �  �  �  �  �  �                             ���   ��������������������Ƅ  �  �  �  �  �  �  �  �  �  �  �  �  �  ������   ������   ������   ���   �����Ƅ�������������Ƅ  �  �  �  �  �  �  �  �  �  �  �  �  �  ������   ������   ������   ���   �����Ƅ����� �������Ƅ  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ���   �����Ƅ�� ����Ƅ�������������������������������������������������������������������������Ƅ��   �����Ƅ��������������������������������������������������������������������������������������   ��������������������������������������������������������������������������Ƅ��   ���������������Ƅ  �  �  �  �  �  �  �  �  �  �  �  �  �                             ���   ���������������Ƅ  �  �  �  �  �  �  �  �  �  �  �  �  �  ������   ������   ������   ���   ���������������Ƅ  �  �  �  �  �  �  �  �  �  �  �  �  �  ������   ������   ������   ���   ���������������Ƅ  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ���   ������������������������������������������������������������������������������������Ƅ��   ����������������������������������������������������������������������������������������   ����������Transparent	OnClickExplorerClick  TRadioButtonCommanderInterfaceButton2LeftTopWidthuHeightCaption
&CommanderChecked	TabOrder TabStop	  TRadioButtonExplorerInterfaceButton2LeftTop� WidthoHeightCaption&UtforskareTabOrder       TPF0TImportSessionsDialogImportSessionsDialogLeftjTop� HelpType	htKeywordHelpKeyword	ui_importBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionImportera sessioner fr�n PuTTYClientHeightClientWidthwColor	clBtnFace
ParentFont	OldCreateOrder	PositionpoMainFormCenterOnClose	FormCloseOnShowFormShow
DesignSizew PixelsPerInch`
TextHeight TLabelLabel1LeftTopWidthiHeight-AnchorsakLeftakTopakRight AutoSizeCaption�F�ljande lista inneh�ller sessioner som har lagrats av SSH-klienten PuTTY. V�lj de sessioner som ska importeras och klicka sedan p� OK.WordWrap	  TButtonOKButtonLeft� Top� WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top� WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  	TListViewSessionListViewLeftTop4WidthiHeight� AnchorsakLeftakTopakRightakBottom 
Checkboxes	ColumnsCaptionSessionWidth�  Caption	ProtokollWidth<  ColumnClickHideSelectionReadOnly	ParentShowHintShowHint	TabOrder 	ViewStylevsReport	OnInfoTipSessionListViewInfoTipOnKeyUpSessionListViewKeyUpOnMouseDownSessionListViewMouseDown  TButtonCheckAllButtonLeftTop� WidthYHeightAnchorsakLeftakBottom CaptionMarkera/avmarkera &allaTabOrderOnClickCheckAllButtonClick  	TCheckBoxImportKeysCheckLeftTop� WidthYHeightAnchorsakLeftakBottom Caption2Importera cachade &v�rdnycklar f�r valda sessionerTabOrder  TButton
HelpButtonLeft&Top� WidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrderOnClickHelpButtonClick     TPF0TLicenseDialogLicenseDialogLeft�Top� ActiveControlCloseButtonBorderIconsbiSystemMenu BorderStylebsDialogCaptionAnv�ndarlicensClientHeight@ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrder	PositionpoMainFormCenter
DesignSize�@ PixelsPerInch`
TextHeight TButtonCloseButtonLeft�TopWidthKHeightAnchorsakRightakBottom Cancel	CaptionSt�ngDefault	ModalResultTabOrder   TMemoLicenseMemoLeftTopWidth�HeightAnchorsakLeftakTopakRight Color	clBtnFaceReadOnly	
ScrollBars
ssVerticalTabOrderWantReturns   TPF0TLocationProfilesDialogLocationProfilesDialogLeftWTop� HelpType	htKeywordHelpKeywordui_locationprofileBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionPlatsprofilerClientHeight�ClientWidth-Color	clBtnFace
ParentFont	OldCreateOrder	PositionpoMainFormCenterOnShowFormShow
DesignSize-� PixelsPerInch`
TextHeight TLabelLocalDirectoryLabelLeftTopWidthHHeightCaptionL&okal katalog:FocusControlLocalDirectoryEdit  TLabelRemoteDirectoryLabelLeftTop8WidthSHeightCaptionF&j�rrkatalog:FocusControlRemoteDirectoryEdit  TButtonOKBtnLeft/Top�WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeft�Top�WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TPageControlPageControlLeftTophWidthHeight 
ActivePageSessionProfilesSheetAnchorsakLeftakTopakRightakBottom TabIndex TabOrder 	TTabSheetSessionProfilesSheetTagCaptionSessionsplatsprofiler
DesignSize  	TTreeViewSessionProfilesViewTagLeft
Top	Width�Height� AnchorsakLeftakTopakRightakBottom DragModedmAutomaticHideSelectionImagesBookmarkImageListIndentTabOrder OnChangeProfilesViewChangeOnCollapsedProfilesViewCollapsed
OnDblClickProfilesViewDblClick
OnDragDropProfilesViewDragDrop
OnDragOverProfilesViewDragOverOnEditedProfilesViewEdited	OnEditingProfilesViewEditing	OnEndDragProfilesViewEndDrag
OnExpandedProfilesViewExpandedOnGetImageIndexProfilesViewGetImageIndexOnGetSelectedIndexProfilesViewGetSelectedIndex	OnKeyDownProfilesViewKeyDownOnStartDragProfilesViewStartDrag
Items.Data
�                ��������       1           ��������        11           ��������        2           ��������        3          ��������       4           ��������        41           ��������        5  TButtonAddSessionBookmarkButtonTagLeft�Top	WidthSHeightAnchorsakTopakRight Caption&L�gg till...TabOrderOnClickAddBookmarkButtonClick  TButtonRemoveSessionBookmarkButtonTagLeft�Top)WidthSHeightAnchorsakTopakRight Caption&Ta bortTabOrderOnClickRemoveBookmarkButtonClick  TButtonDownSessionBookmarkButtonTagLeft�Top� WidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickBookmarkButtonClick  TButtonUpSessionBookmarkButtonTag�Left�Top� WidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickBookmarkButtonClick  TButtonRenameSessionBookmarkButtonTagLeft�TopIWidthSHeightAnchorsakTopakRight Caption	B&yt namnTabOrderOnClickRenameBookmarkButtonClick  TButtonSessionBookmarkMoveToButtonTagLeft�TopiWidthSHeightAnchorsakTopakRight Caption&Flytta till...TabOrderOnClickBookmarkMoveToButtonClick   	TTabSheetSharedProfilesSheetTagCaptionDelade platsprofiler
ImageIndex
DesignSize  	TTreeViewSharedProfilesViewTagLeft
Top	Width�Height� AnchorsakLeftakTopakRightakBottom DragModedmAutomaticHideSelectionImagesBookmarkImageListIndentTabOrder OnChangeProfilesViewChangeOnCollapsedProfilesViewCollapsed
OnDblClickProfilesViewDblClick
OnDragDropProfilesViewDragDrop
OnDragOverProfilesViewDragOverOnEditedProfilesViewEdited	OnEditingProfilesViewEditing	OnEndDragProfilesViewEndDrag
OnExpandedProfilesViewExpandedOnGetImageIndexProfilesViewGetImageIndexOnGetSelectedIndexProfilesViewGetSelectedIndex	OnKeyDownProfilesViewKeyDownOnStartDragProfilesViewStartDrag
Items.Data
�                ��������       1           ��������        11           ��������        2           ��������        3          ��������       4           ��������        41           ��������        5  TButtonAddSharedBookmarkButtonTagLeft�Top	WidthSHeightAnchorsakTopakRight Caption&L�gg till...TabOrderOnClickAddBookmarkButtonClick  TButtonRemoveSharedBookmarkButtonTagLeft�Top)WidthSHeightAnchorsakTopakRight Caption&Ta bortTabOrderOnClickRemoveBookmarkButtonClick  TButtonRenameSharedBookmarkButtonTagLeft�TopIWidthSHeightAnchorsakTopakRight Caption	B&yt namnTabOrderOnClickRenameBookmarkButtonClick  TButtonSharedBookmarkMoveToButtonTagLeft�TopiWidthSHeightAnchorsakTopakRight Caption&Flytta till...TabOrderOnClickBookmarkMoveToButtonClick  TButtonUpSharedBookmarkButtonTag�Left�Top� WidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickBookmarkButtonClick  TButtonDownSharedBookmarkButtonTagLeft�Top� WidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickBookmarkButtonClick  TButtonShortCutSharedBookmarkButtonTagLeft�Top� WidthSHeightAnchorsakTopakRight Caption
&Genv�g...TabOrderOnClickShortCutBookmarkButtonClick    TIEComboBoxLocalDirectoryEditLeftTopWidth�HeightAnchorsakLeftakTopakRight 
ItemHeightTabOrder TextLocalDirectoryEditOnChangeDirectoryEditChange  TIEComboBoxRemoteDirectoryEditLeftTopIWidthHeightAnchorsakLeftakTopakRight 
ItemHeight	MaxLength�TabOrderTextRemoteDirectoryEditOnChangeDirectoryEditChange  TButtonLocalDirectoryBrowseButtonLeft�TopWidthKHeightAnchorsakTopakRight CaptionBl�dd&ra...TabOrderOnClickLocalDirectoryBrowseButtonClick  TButtonSwitchButtonLeftTop�WidthaHeightAnchorsakRightakBottom Caption&Bokm�rken...ModalResultTabOrderOnClickSwitchButtonClick  TButton
HelpButtonLeft�Top�WidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrderOnClickHelpButtonClick  
TImageListBookmarkImageListLeft� Top�Bitmap
&  IL     �������������BM6       6   (   @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            !! !! !! !! !! !! !! !! !! !! !! !! !!                                                                                         ff ���  ��  ��  ��  ��  ��  ��  ��  ��  ��  �� f��  ��              ff  ff  ff  ff  ff  ff  ff  ff  ff  ff  ff  ff !! !!      ff ���  ��  ��  ��  ��  ��  ��  ��  ��  �� f��  �� f��                                                                       ff ���  ��  ��  ��  ��  �� �    ��  ��  ��  ��  �� f��              ff ���  ��  ��  ��  ��  ��  ��  �� f��  ��  ff !! !!      ff ���  ��  ��  ��  ��  ��  ��  ��  ��  ��  �� f��  ��                                                                       ff ��� ���  ��  �� �    �� �    �� �    ��  ��  ��  ��          ff ���  ��  ��  ��  ��  ��  ��  ��  ��  �� f�� !!  ff !!      ff ��� ���  ��  ��  ��  ��  ��  ��  ��  ��  ��  �� f��                                                                       ff ���  �� ���  ��  �� �   �   �    ��  ��  ��  ��  ��          ff ��� ���  ��  ��  ��  ��  ��  ��  ��  ��  �� !!  ff !!      ff ���  �� ���  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��                                                                       ff ��� ���  �� �   �   �    �� �   �   �    ��  ��  ��      ff ��� ���  �� ���  ��  ��  ��  ��  ��  ��  �� !!  ��  �� !!      ff ��� ���  �� ���  ��  ��  ��  ��  ��  ��  ��  ��  ��                                                                       ff ���  �� ���  ��  �� �   �   �    ��  ��  ��  ��  ��      ff ���  �� ���  �� ���  ��  ��  ��  ��  ��  �� !!  ��  �� !!      ff ���  �� ���  �� ���  �� ���  ��  ��  ��  ��  ��  ��                                                                       ff ��� ���  �� ��� �    �� �    �� �    ��  ��  ��  ��      ff  ff  ff  ff  ff  ff  ff  ff  ff  ff  ff  ff  ��  ��  �� !!      ff ��� ���  �� ���  �� ���  �� ���  ��  ��  ��  ��  ��                                                                       ff ���  �� ���  �� ���  �� �    ��  ��  ��  ��  ��  ��          ff ���  �� ���  ��  ��  ��  ��  ��  ��  ��  ��  ��  �� !!      ff ���  �� ���  �� ���  �� ���  �� ���  ��  ��  ��  ��                                                                       ff ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���          ff ��� ���  �� ���  ��  ��  ��  �� ��� ��� ��� ��� ��� !!      ff ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                       ff  ff  ff  ff  ff  ff  ff  ff  ff  ff  ff  ff  ff  ff          ff ���  �� ���  �� ���  �� ���  ff  ff  ff  ff  ff  ff          ff  ff  ff  ff  ff  ff  ff  ff  ff  ff  ff  ff  ff  ff                                                                           ff ��� ��� ��� ��� ���                                          ff ��� ��� ��� ��� ���  ff                                      ff ��� ��� ��� ���  ��                                                                                                           ff  ff  ff  ff  ff                                              ff  ff  ff  ff  ff                                              ff  ff  ff  ff  ff                                                                                                                                                                                                                                                                                                                                                                 BM>       >   (   @            �                       ��� ������  ������  � � �   � � �   � � �   � � �   � � �   �   �   �   �   �   �   � � �   � � �   � ��   ���  ������  ������                           TPF0TLogFormLogFormLeftdTop� Width�HeightUHelpType	htKeywordHelpKeywordui_logBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp CaptionLogColor	clBtnFaceConstraints.MinHeight� Constraints.MinWidth� Font.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameMS Sans Serif
Font.Style 	Icon.Data
6           (  &          �  N  (                �                         �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���          33330  �����  �����  �����  ����  ��w��  ���  �����  ���x�  �����  �����  ���x�  �����  �����         ��  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  (       @         �                        �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                                   33333333330     ����������     �����������     o���������     ���������     �����������     o�����x���     ���������     ���������     o���������     ����xx��     ��������     o���8����     ���?������     �����������     o����������     ���8���Ǐ�     ����?��̏��     o���8���x��     ���?��̏��     ����8���x��     o���?��̏��     �������x��     �������̏��     o����������     ����������     �����������                                                  �����  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ��������OldCreateOrderPositionpoDefaultPosOnlyOnClose	FormClosePixelsPerInch`
TextHeight TTBXStatusBar	StatusBarLeft Top Width�HeightPanelsFramedMaxSize� Size� StretchPrioritydTag   UseSystemFont  TTBXDockTopDockLeft Top Width�Height	AllowDrag TTBXToolbarToolbarLeft Top CaptionToolbarFullSize	ImagesGlyphsModule.LogImagesParentShowHintShowHint	TabOrder  TTBXItemTBXItem1Action"NonVisualDataModule.LogCloseAction  TTBXSeparatorItemTBXSeparatorItem1  TTBXItemTBXItem2Action"NonVisualDataModule.LogClearAction  TTBXItemTBXItem3Action!NonVisualDataModule.LogCopyAction  TTBXItemTBXItem4Action&NonVisualDataModule.LogSelectAllAction  TTBXSeparatorItemTBXSeparatorItem2  TTBXItemTBXItem5Action(NonVisualDataModule.LogPreferencesAction        TPF0TLoggingFrameLoggingFrameLeft Top Width:HeightTabOrder 
DesignSize:  	TGroupBoxLoggingGroupLeftTop;Width5Height� AnchorsakLeftakTopakRight CaptionAlternativ f�r loggningTabOrder 
DesignSize5�   TLabelLogWindowLinesTextLeft Top� WidthHeightCaptionrader  TLabelLogProtocolLabelLeftTopWidthBHeightCaptionNiv� &loggning:FocusControlLogProtocolCombo  	TCheckBoxLogToFileCheckLeftTop-Width� HeightCaptionLogga till &fil:TabOrderOnClickLogToFileCheckChange  TFilenameEditLogFileNameEdit2Left(TopDWidth� HeightAcceptFiles	OnBeforeDialogLogFileNameEdit2BeforeDialogOnAfterDialogLogFileNameEdit2AfterDialog
DefaultExtlogFilter9Loggfiler (*.log; *.xml)|*.log;*.xml|Alla filer (*.*)|*.*DialogOptionsofHideReadOnlyofPathMustExist DialogTitleV�lj fil f�r sessionsloggen.OnCreateEditDialog LogFileNameEdit2CreateEditDialogClickKey@AnchorsakLeftakTopakRight TabOrderTextLogFileNameEdit2OnChange
DataChange  	TCheckBoxLogShowWindowCheckLeftTopyWidth� HeightCaptionVisa loggf&�nster:TabOrderOnClick
DataChange  TRadioButtonLogWindowCompleteButtonLeft(Top� Width� HeightCaptionVisa &hela sessionenTabOrderOnClick
DataChange  TRadioButtonLogWindowLinesButtonLeft(Top� Width� HeightCaptionVisa endast &senasteTabOrderOnClick
DataChange  TUpDownEditLogWindowLinesEditLeft� Top� WidthIHeight	AlignmenttaRightJustify	Increment2MaxValue'MinValue2Value2TabOrderOnChange
DataChange  TPanelLogFilePanelLeft(Top]Width� HeightAnchorsakLeftakTopakRight 
BevelOuterbvNoneTabOrder TRadioButtonLogFileAppendButtonLeft TopWidthaHeightCaption
L&�gg tillTabOrder OnClick
DataChange  TRadioButtonLogFileOverwriteButtonLeft`TopWidthYHeightCaptionSk&riv �verTabOrderOnClick
DataChange   	TComboBoxLogProtocolComboLeftpTopWidthqHeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrder Items.StringsNormalDebug 1Debug 2   TStaticTextLogFileNameHintTextLeft� Top[WidthGHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption&m�nsterTabOrderTabStop	   	TGroupBoxLogGroupLeftTopWidth5Height3AnchorsakLeftakTopakRight CaptionLoggTabOrder TRadioButtonLoggingOffButtonLeftTopWidthYHeightCaptionI&ngen loggTabOrder OnClickLoggingButtonClick  TRadioButtonLoggingOnButtonLeftpTopWidthYHeightCaption
&Text loggTabOrderOnClickLoggingButtonClick  TRadioButtonLoggingActionsButtonLeft� TopWidthYHeightCaption	&XML loggTabOrderOnClickLoggingButtonClick     TPF0TLoginDialogLoginDialogLeft_Top� HelpType	htKeywordHelpKeywordui_loginBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption
InloggningClientHeightPClientWidthColor	clBtnFace
ParentFont	
KeyPreview	OldCreateOrder	PositionpoMainFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSizeP PixelsPerInch`
TextHeight TButton
HelpButtonLeft�Top1WidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrderVisibleOnClickHelpButtonClick  TButton
SaveButtonLeftSTop1WidthKHeightHelpKeywordui_login_saveActionSaveSessionActionAnchorsakRightakBottom TabOrder  TButtonLoginButtonLeft� Top1WidthKHeightActionLoginActionAnchorsakRightakBottom Default	ModalResultTabOrder  TButtonCloseButtonLeft�Top1WidthKHeightAnchorsakRightakBottom Cancel	CaptionSt�ngModalResultTabOrder  TButtonAboutButtonLeftTop1WidthRHeightActionAboutActionAnchorsakLeftakBottom TabOrder TabStop  TButtonLanguagesButtonLeftiTop1WidthKHeightAnchorsakLeftakBottom Caption
Lan&guagesTabOrderOnClickLanguagesButtonClick  TPanel	MainPanelLeft Top WidthHeight(AlignalTopAnchorsakLeftakTopakRightakBottom 
BevelOuterbvNoneTabOrder TPageControlPageControlTagLeft� Top WidthiHeight(HelpType	htKeyword
ActivePage
BasicSheetAlignalClient	MultiLine	Style	tsButtonsTabOrderTabStopOnChangePageControlChange 	TTabSheet
BasicSheetTagHintSessionHelpType	htKeywordHelpKeywordui_login_sessionCaptionBasic
ImageIndex
TabVisible
DesignSizea  	TGroupBox
BasicGroupLeft TopWidthYHeight� AnchorsakLeftakTopakRight CaptionSessionTabOrder 
DesignSizeY�   TLabelLabel1LeftTopWidth6HeightCaption
&V�rdnamn:FocusControlHostNameEdit  TLabelLabel2Left� TopWidth<HeightAnchorsakTopakRight CaptionPo&rtnummer:FocusControlPortNumberEdit  TLabelLabel3LeftTopDWidth6HeightCaption&Anv�ndarnamn:FocusControlUserNameEdit  TLabelLabel4Left� TopDWidth1HeightCaption
&L�senord:FocusControlPasswordEdit  TLabelPrivateKeyLabelLeftTopvWidthHHeightCaptionFil med privat nyc&kelFocusControlPrivateKeyEdit  TEditHostNameEditLeftTop#Width� HeightAnchorsakLeftakTopakRight 	MaxLengthdTabOrder TextHostNameEditOnChange
DataChange  TEditUserNameEditLeftTopUWidth� Height	MaxLengthdTabOrderTextUserNameEditOnChange
DataChange  TPasswordEditPasswordEditLeft� TopUWidth� HeightAnchorsakLeftakTopakRight 	MaxLengthdTabOrderTextPasswordEditOnChange
DataChange  TUpDownEditPortNumberEditLeft� Top#WidthRHeight	AlignmenttaRightJustifyMaxValue��  MinValueValueAnchorsakTopakRight TabOrderOnChange
DataChange  TFilenameEditPrivateKeyEditLeftTop� WidthBHeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPrivateKeyEditAfterDialogFilter8PuTTY privata nycklar (*.ppk)|*.ppk|Alla filer (*.*)|*.*DialogOptions
ofReadOnlyofPathMustExistofFileMustExist DialogTitleV�lj privat nyckelfilClickKey@AnchorsakLeftakTopakRight TabOrderTextPrivateKeyEditOnChange
DataChange   	TGroupBoxTransferProtocolGroupLeft Top� WidthYHeight/AnchorsakLeftakTopakRight Caption	ProtokollTabOrder TLabelLabel22LeftTopWidth<HeightCaption&Filprotokoll:FocusControlTransferProtocolCombo  	TComboBoxTransferProtocolComboLeftlTopWidth;HeightStylecsDropDownList
ItemHeightTabOrder OnChangeTransferProtocolComboChangeItems.StringsSFTPSCPFTP   	TCheckBoxAllowScpFallbackCheckLeft� TopWidthyHeightCaptionTill�t SCP &fallbackTabOrderOnClick
DataChange  	TComboBox	FtpsComboLeft� TopWidth� HeightStylecsDropDownList
ItemHeightTabOrderOnChangeTransferProtocolComboChangeItems.StringsIngen krypteringSSL/TLS Implicit encryptionXSSL Explicit encryptionXTLS Explicit encryptionX    TButtonColorButtonLeftTop� WidthKHeightCaption
V�lj f&�rgTabOrderOnClickColorButtonClick   	TTabSheetSessionListSheetTagHintLagrade sessionerHelpType	htKeywordHelpKeywordui_login_stored_sessionsCaptionStSe
TabVisible
DesignSizea  TButton
LoadButtonLeftTop#WidthXHeightActionEditSessionActionAnchorsakTopakRight TabOrder  TButtonDeleteButtonLeftTopCWidthXHeightActionDeleteSessionActionAnchorsakTopakRight TabOrder  	TTreeViewSessionTreeLeftTopWidth� HeightAnchorsakLeftakTopakRightakBottom DragModedmAutomaticHideSelectionIndentParentShowHint	RowSelect	ShowHint		ShowLinesShowRootSortTypestBothStateImagesSessionImageListTabOrder OnChangeSessionTreeChangeOnCollapsedSessionTreeExpandedCollapsed	OnCompareSessionTreeCompareOnCustomDrawItemSessionTreeCustomDrawItem
OnDblClickSessionTreeDblClick
OnDragDropSessionTreeDragDropOnEditedSessionTreeEdited	OnEditingSessionTreeEditing	OnEndDragSessionTreeEndDrag
OnExpandedSessionTreeExpandedCollapsed	OnKeyDownSessionTreeKeyDownOnMouseMoveSessionTreeMouseMoveOnStartDragSessionTreeStartDrag  TButton	NewButtonLeftTopWidthXHeightActionNewSessionActionAnchorsakTopakRight TabOrder  TButtonSetDefaultSessionButtonLeftTop� WidthXHeightActionSetDefaultSessionActionAnchorsakTopakRight TabOrder  TButtonToolsMenuButtonLeftTopWidthXHeightAnchorsakRightakBottom Caption&Verktyg...TabOrderOnClickToolsMenuButtonClick  TButtonShellIconsButtonLeftTop� WidthXHeightActionShellIconSessionActionAnchorsakTopakRight TabOrder  TButtonRenameButtonLeftTopcWidthXHeightActionRenameSessionActionAnchorsakTopakRight TabOrder  TButtonNewFolderButtonLeftTop� WidthXHeightActionNewSessionFolderActionAnchorsakTopakRight TabOrder   	TTabSheetLogSheetTagHintLoggningHelpType	htKeywordHelpKeywordui_login_loggingCaptionLog
ImageIndex
TabVisible �TLoggingFrameLoggingFrameLeft�Top WidthdHeightTabOrder 
DesignSized  �	TGroupBoxLoggingGroupWidthY �	TCheckBoxLogToFileCheckWidth9  �TFilenameEditLogFileNameEdit2Width#  �	TCheckBoxLogShowWindowCheckWidthA  �TRadioButtonLogWindowCompleteButtonWidth!  �TPanelLogFilePanelWidth# �TRadioButtonLogFileAppendButtonCaption
&L�gg till  �TRadioButtonLogFileOverwriteButtonWidth�    �TStaticTextLogFileNameHintTextLeft    �	TGroupBoxLogGroupWidthY    	TTabSheetEnvironmentSheetTagHintMilj�HelpType	htKeywordHelpKeywordui_login_environmentCaptionEnv
ImageIndex
TabVisible
DesignSizea  TLabelEnvironmentOtherLabelLeft Top� WidthDHeightCaption�vriga inst�llningar:  TStaticTextRecycleBinLinkLabelLeftXTop� Width<HeightCaptionPapperskorgTabOrderTabStop	OnClickRecycleBinLinkLabelClick  	TGroupBoxEnvironmentGroupLeft TopWidthYHeight`AnchorsakLeftakTopakRight CaptionServermilj�TabOrder 
DesignSizeY`  TLabelEOLTypeLabelLeftTopWidth� HeightCaption0Slut p� rad &tecken (om det inte ges av server):FocusControlEOLTypeCombo  TLabelUtfLabelLeftTop,Width� HeightCaption&UTF-8 kodning p� filnamn:FocusControlUtfCombo  TLabelTimeDifferenceLabelLeftTopDWidthNHeightCaptionOffset tidszon:FocusControlTimeDifferenceEdit  TLabelTimeDifferenceHoursLabelLeft� TopDWidthHeightCaptiontimmarFocusControlTimeDifferenceEdit  TLabelTimeDifferenceMinutesLabelLeft(TopBWidth$HeightCaptionminuterFocusControlTimeDifferenceMinutesEdit  	TComboBoxEOLTypeComboLeftTopWidth=HeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrder Items.StringsLFCR/LF   	TComboBoxUtfComboLeftTop'Width=HeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrder  TUpDownEditTimeDifferenceEditLeft� Top?Width6Height	AlignmenttaRightJustifyMaxValueMinValue�Value�AnchorsakTopakRight TabOrderOnChange
DataChange  TUpDownEditTimeDifferenceMinutesEditLeft� Top?Width6Height	AlignmenttaRightJustify	IncrementMaxValue-MinValue�Value�AnchorsakTopakRight TabOrderOnChange
DataChange   	TGroupBoxDSTModeGroupLeft TopnWidthYHeight]AnchorsakLeftakTopakRight Caption	SommartidTabOrder
DesignSizeY]  TRadioButtonDSTModeUnixCheckLeftTopWidth=HeightAnchorsakLeftakTopakRight Caption5Justera fj�rrtidsst�mpel med lokal ko&nvention (Unix)TabOrder OnClick
DataChange  TRadioButtonDSTModeWinCheckLeftTop*Width=HeightAnchorsakLeftakTopakRight Caption+Justera fj�rrtidsst�mpel med &DST (Windows)TabOrderOnClick
DataChange  TRadioButtonDSTModeKeepCheckLeftTopAWidth=HeightAnchorsakLeftakTopakRight CaptionBevara fj�rrtidsst�mpel (Unix)TabOrderOnClick
DataChange    	TTabSheetDirectoriesSheetTagHint	KatalogerHelpType	htKeywordHelpKeywordui_login_directoriesCaptionDir
ImageIndex
TabVisible
DesignSizea  	TGroupBoxDirectoriesGroupLeft TopWidthYHeight� AnchorsakLeftakTopakRight Caption	KatalogerTabOrder 
DesignSizeY�   TLabelLocalDirectoryLabelLeftTopTWidthHHeightCaption&Lokal katalogFocusControlLocalDirectoryEdit  TLabelRemoteDirectoryLabelLeftTop)WidthSHeightCaptionF&j�rrkatalogFocusControlRemoteDirectoryEdit  TLabelLocalDirectoryDescLabelLeftTop~Width� HeightCaption@Lokal katalog anv�nds inte i det utforskar-liknande gr�nssnittet  TDirectoryEditLocalDirectoryEditLeftTopeWidthCHeightAcceptFiles	
DialogTextV�lj lokal katalog vid uppstartClickKey@AnchorsakLeftakTopakRight TabOrderTextLocalDirectoryEditOnChange
DataChange  TEditRemoteDirectoryEditLeftTop:WidthCHeightAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextRemoteDirectoryEditOnChange
DataChange  	TCheckBoxUpdateDirectoriesCheckLeftTopWidthAHeightAnchorsakLeftakTopakRight Caption Ko&m ih�g senast anv�nda katalogTabOrder    	TGroupBoxDirectoryOptionsGroupLeft Top� WidthYHeightWAnchorsakLeftakTopakRight CaptionAlternativ vid kalalogl�sningTabOrder
DesignSizeYW  	TCheckBoxCacheDirectoriesCheckLeftTopWidthAHeightAnchorsakLeftakTopakRight CaptionCacha &bes�kta fj�rrkatalogerTabOrder OnClick
DataChange  	TCheckBoxCacheDirectoryChangesCheckLeftTop'Width� HeightAnchorsakLeftakTopakRight CaptionCacha katalogf&�r�ndringarTabOrderOnClick
DataChange  	TCheckBoxResolveSymlinksCheckLeftTop;WidthAHeightAnchorsakLeftakTopakRight CaptionSl� upp symboliska l�&nkarTabOrder  	TCheckBoxPreserveDirectoryChangesCheckLeft� Top'Width� HeightAnchorsakLeftakTopakRight Caption&Permanent cacheTabOrder    	TTabSheetRecycleBinSheetTagHintPapperskorgHelpType	htKeywordHelpKeywordui_login_recycle_binCaptionRec
ImageIndex
TabVisible
DesignSizea  	TGroupBoxRecycleBinGroupLeft TopWidthYHeightrAnchorsakLeftakTopakRight CaptionPapperskorgTabOrder 
DesignSizeYr  TLabelRecycleBinPathLabelLeftTop@Width^HeightCaptionPapp&erskorg p� servernFocusControlRecycleBinPathEdit  	TCheckBoxDeleteToRecycleBinCheckLeftTopWidth=HeightCaption5Flytta borttagna filer p� servern till &papperskorgenTabOrder OnClick
DataChange  	TCheckBoxOverwrittenToRecycleBinCheckLeftTop*Width=HeightCaptionEFlytta &�verskrivna filer p� servern till papperskorgen (endast SFTP)TabOrderOnClick
DataChange  TEditRecycleBinPathEditLeftTopQWidthBHeightAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextRecycleBinPathEditOnChange
DataChange    	TTabSheet	SftpSheetTagHintSFTPHelpType	htKeywordHelpKeywordui_login_sftpCaptionSftp
ImageIndex
TabVisible
DesignSizea  	TGroupBoxSFTPBugsGroupBoxLeft TopTWidthYHeightFAnchorsakLeftakTopakRight CaptionUppt�ckta buggar i SFTP servrarTabOrder
DesignSizeYF  TLabelLabel10LeftTopWidth� HeightCaption8&Omv�nd ordning p� symboliska l�nkar i kommandoargument:FocusControlSFTPBugSymlinkCombo  TLabelLabel36LeftTop,Width� HeightCaption1Feltolkning av filtidsst�&mplar tidigare �n 1970:FocusControlSFTPBugSignedTSCombo  	TComboBoxSFTPBugSymlinkComboLeftTopWidth=HeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrder   	TComboBoxSFTPBugSignedTSComboLeftTop'Width=HeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrder   	TGroupBoxSFTPProtocolGroupLeft TopWidthYHeightFAnchorsakLeftakTopakRight CaptionAlternativ f�r protokollTabOrder 
DesignSizeYF  TLabelLabel34LeftTop,Width� HeightCaption!F�re&drar SFTP protokoll version:FocusControlSFTPMaxVersionCombo  TLabelLabel23LeftTopWidth>HeightCaptionSFTP ser&verFocusControlSftpServerEdit  	TComboBoxSFTPMaxVersionComboLeftTop'Width=HeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrderItems.Strings012345   	TComboBoxSftpServerEditLeft� TopWidth� HeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeight	MaxLength� TabOrder TextSftpServerEditItems.StringsStandard/bin/sftp-serversudo su -c /bin/sftp-server     	TTabSheetScpSheetTagHintSCP/SkalHelpType	htKeywordHelpKeywordui_login_scpCaptionShl
ImageIndex
TabVisible
DesignSizea  	TGroupBoxOtherShellOptionsGroupLeft Top� WidthYHeightEAnchorsakLeftakTopakRight Caption�vriga alternativTabOrder 	TCheckBoxLookupUserGroupsCheckLeftTopWidth� HeightCaptionSl� upp &anv�ndargrupperTabOrder OnClick
DataChange  	TCheckBoxClearAliasesCheckLeftTop*Width� HeightCaptionRensa a&liasTabOrderOnClick
DataChange  	TCheckBoxUnsetNationalVarsCheckLeft� TopWidth� HeightCaptionRensa &nationella variablerTabOrderOnClick
DataChange  	TCheckBoxScp1CompatibilityCheckLeft� Top*Width� HeightCaption$Anv�nd scp&2 med scp1 kompatibilitetTabOrderOnClick
DataChange   	TGroupBox
ShellGroupLeft TopWidthYHeightFAnchorsakLeftakTopakRight CaptionSkalTabOrder 
DesignSizeYF  TLabelLabel19LeftTopWidthHeightCaptionS&kal:FocusControl	ShellEdit  TLabelLabel20LeftTop,WidthfHeightCaption&Returnera kodvariabel:FocusControlReturnVarEdit  	TComboBox	ShellEditLeft� TopWidth� HeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeight	MaxLength2TabOrder Text	ShellEditItems.StringsStandard	/bin/bash/bin/ksh	sudo su -   	TComboBoxReturnVarEditLeft� Top'Width� HeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeight	MaxLength2TabOrderTextReturnVarEditItems.StringsDetektera automatiskt?status    	TGroupBoxScpLsOptionsGroupLeft TopTWidthYHeightEAnchorsakLeftakTopakRight CaptionListning av katalogerTabOrder
DesignSizeYE  TLabelLabel9LeftTopWidthRHeightCaption&Kommando f�r listning:FocusControlListingCommandEdit  	TCheckBoxIgnoreLsWarningsCheckLeftTop*Width� HeightCaptionIgnorera LS &varningarTabOrderOnClick
DataChange  	TCheckBoxSCPLsFullTimeAutoCheckLeft� Top*Width� HeightCaptionF�rs�k att f� &full tidsst�mpelTabOrderOnClick
DataChange  	TComboBoxListingCommandEditLeft� TopWidth� HeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeight	MaxLength2TabOrder TextListingCommandEditItems.Stringsls -lals -gla     	TTabSheetFtpSheetTagHintFTPHelpType	htKeywordHelpKeywordui_login_ftpCaptionFtpSheet
ImageIndex
TabVisible
DesignSizea  	TGroupBoxFtpGroupLeft TopWidthYHeight� AnchorsakLeftakTopakRight CaptionAlternativ f�r protokollTabOrder 
DesignSizeY�   TLabelLabel25LeftTopWidthgHeightCaption&Kommandon efter inloggning:FocusControlPostLoginCommandsMemo  TLabelLabel5LeftTopfWidth� HeightCaption$&Support f�r listning av dolda filerFocusControlFtpListAllCombo  TMemoPostLoginCommandsMemoLeftTop%WidthAHeight5AnchorsakLeftakTopakRight 	MaxLength2
ScrollBars
ssVerticalTabOrder   	TComboBoxFtpListAllComboLeftTopaWidth=HeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrder  	TCheckBoxFtpForcePasvIpCheckLeftTop}Width=HeightCaption*&Tvinga ip-adress f�r passiva anslutningarTabOrderOnClick
DataChange    	TTabSheet	ConnSheetTagHint
AnslutningHelpType	htKeywordHelpKeywordui_login_connectionCaptionConn
ImageIndex
TabVisible
DesignSizea  	TGroupBoxFtpPingGroupLeft ToplWidthYHeightuAnchorsakLeftakTopakRight Caption
KeepalivesTabOrder
DesignSizeYu  TLabelFtpPingIntervalLabelLeftTopZWidth� HeightCaptionSekunder &mellan keepalivesFocusControlFtpPingIntervalSecEdit  TUpDownEditFtpPingIntervalSecEditLeft� TopUWidthIHeight	AlignmenttaRightJustifyMaxValueMinValue	MaxLengthTabOrderOnChange
DataChange  TRadioButtonFtpPingOffButtonLeftTopWidth=HeightAnchorsakLeftakTopakRight Caption&AvTabOrder OnClick
DataChange  TRadioButtonFtpPingNullPacketButtonLeftTop*Width=HeightAnchorsakLeftakTopakRight CaptionSkicka SSH-&null-paketEnabledTabOrderOnClick
DataChange  TRadioButtonFtpPingDummyCommandButtonLeftTopAWidth=HeightAnchorsakLeftakTopakRight Caption!K�r kommandon f�r &dummy-protkollTabOrderOnClick
DataChange   	TGroupBoxTimeoutGroupLeft Top9WidthYHeight.AnchorsakLeftakTopakRight Caption	TimeouterTabOrder TLabelLabel11LeftTopWidthuHeightCaptionTimeout f�r se&rversvar:FocusControlTimeoutEdit  TLabelLabel12LeftTopWidth(HeightCaptionsekunderFocusControlTimeoutEdit  TUpDownEditTimeoutEditLeft� TopWidthIHeight	AlignmenttaRightJustify	IncrementMaxValuepMinValue	MaxLengthTabOrder OnChange
DataChange   	TGroupBox	PingGroupLeft ToplWidthYHeightuAnchorsakLeftakTopakRight Caption
KeepalivesTabOrder
DesignSizeYu  TLabelPingIntervalLabelLeftTopZWidth� HeightCaptionSekunder &mellan keepalivesFocusControlPingIntervalSecEdit  TUpDownEditPingIntervalSecEditLeft� TopUWidthIHeight	AlignmenttaRightJustifyMaxValueMinValue	MaxLengthTabOrderOnChange
DataChange  TRadioButtonPingOffButtonLeftTopWidth=HeightAnchorsakLeftakTopakRight CaptionA&vTabOrder OnClick
DataChange  TRadioButtonPingNullPacketButtonLeftTop*Width=HeightAnchorsakLeftakTopakRight CaptionSkicka SSH-&null-paketTabOrderOnClick
DataChange  TRadioButtonPingDummyCommandButtonLeftTopAWidth=HeightAnchorsakLeftakTopakRight Caption#K�r kommandon f�r &dummy-protokoll:TabOrderOnClick
DataChange   	TGroupBoxIPvGroupLeft Top� WidthYHeight.AnchorsakLeftakTopakRight CaptionVersion f�r internetprotokollTabOrder
DesignSizeY.  TRadioButtonIPAutoButtonLeftTopWidtheHeightAnchorsakLeftakTopakRight CaptionA&utomatiskTabOrder OnClick
DataChange  TRadioButton
IPv4ButtonLeft|TopWidtheHeightAnchorsakLeftakTopakRight CaptionIPv&4TabOrderOnClick
DataChange  TRadioButton
IPv6ButtonLeft� TopWidtheHeightAnchorsakLeftakTopakRight CaptionIPv&6TabOrderOnClick
DataChange   	TGroupBoxConnectionGroupLeft TopWidthYHeight.AnchorsakLeftakTopakRight Caption
AnslutningTabOrder 
DesignSizeY.  	TCheckBoxFtpPasvModeCheckLeftTopWidthAHeightAnchorsakLeftakTopakRight Caption&Passivt l�geTabOrder OnClick
DataChange    	TTabSheet
ProxySheetTagHintProxyHelpType	htKeywordHelpKeywordui_login_proxyCaptionProxy
ImageIndex
TabVisible
DesignSizea  	TGroupBoxProxyTypeGroupLeft TopWidthYHeight� AnchorsakLeftakTopakRight CaptionProxyTabOrder 
DesignSizeY�   TLabelProxyMethodLabelLeftTopWidth4HeightCaption&Typ av proxy:FocusControlSshProxyMethodCombo  TLabelProxyHostLabelLeftTop)WidthQHeightCaptionPro&xyns v�rdnamn:FocusControlProxyHostEdit  TLabelProxyPortLabelLeft� Top)Width<HeightAnchorsakTopakRight CaptionPo&rtnummer:FocusControlProxyPortEdit  TLabelProxyUsernameLabelLeftTopUWidth6HeightCaption&Anv�ndarnamn:FocusControlProxyUsernameEdit  TLabelProxyPasswordLabelLeft� TopUWidth1HeightCaption
&L�senord:FocusControlProxyPasswordEdit  	TComboBoxSshProxyMethodComboLeft� TopWidthnHeightStylecsDropDownList
ItemHeightTabOrder OnChange
DataChangeItems.StringsIngenSOCKS4SOCKS5HTTPTelnetLokal   TUpDownEditProxyPortEditLeft� Top:WidthRHeight	AlignmenttaRightJustifyMaxValue��  MinValueValueAnchorsakTopakRight TabOrderOnChange
DataChange  TEditProxyHostEditLeftTop:Width� HeightAnchorsakLeftakTopakRight 	MaxLength2TabOrderTextProxyHostEditOnChange
DataChange  TEditProxyUsernameEditLeftTopfWidth� Height	MaxLength2TabOrderTextProxyUsernameEditOnChange
DataChange  TPasswordEditProxyPasswordEditLeft� TopfWidth� HeightAnchorsakLeftakTopakRight 	MaxLength2TabOrderTextProxyPasswordEditOnChange
DataChange  	TComboBoxFtpProxyMethodComboLeft� TopWidth� HeightStylecsDropDownListDropDownCount
ItemHeightTabOrderOnChange
DataChangeItems.StringsIngenSOCKS4SOCKS5HTTP
SITE %host!USER %proxyuser, USER %user@%host
OPEN %hostUSER %proxyuser, USER %userUSER %user@%hostUSER %proxyuser@%hostUSER %user@%host %proxyuserUSER %user@%proxyuser@%host    	TGroupBoxProxySettingsGroupLeft Top� WidthYHeight� AnchorsakLeftakTopakRight CaptionInst�llningar proxyTabOrder
DesignSizeY�   TLabelProxyTelnetCommandLabelLeftTopWidthRHeightCaptionTelnetko&mmando:FocusControlProxyTelnetCommandEdit  TLabelLabel17LeftTopcWidth� HeightCaption+L�t &DNS-namnuppslagningar g�ras av proxyn:  TLabelProxyLocalCommandLabelLeftTopWidthjHeightCaptionLokalt proxyko&mmando:FocusControlProxyLocalCommandEdit  TEditProxyTelnetCommandEditLeftTop#WidthBHeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder TextProxyTelnetCommandEditOnChange
DataChange  	TCheckBoxProxyLocalhostCheckLeftTopMWidth9HeightCaption&L�t lokala a&nslutningar g� via proxynTabOrder  	TComboBoxProxyDNSComboLeft� Top^WidthRHeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrderItems.Strings
AutomatiskNejJa   TEditProxyLocalCommandEditLeftTop#Width� HeightAnchorsakLeftakTopakRight TabOrderTextProxyLocalCommandEditOnChange
DataChange  TButtonProxyLocalCommandBrowseButtonLeft� Top!WidthRHeightAnchorsakTopakRight Caption&Bl�ddra...TabOrderOnClick"ProxyLocalCommandBrowseButtonClick  TStaticTextProxyTelnetCommandHintTextLeft� Top:WidthOHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaptionm�nsterTabOrderTabStop	  TStaticTextProxyLocalCommandHintTextLeft� Top:WidthOHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaptionm�nsterTabOrderTabStop	    	TTabSheetTunnelSheetTagHintTunnelHelpType	htKeywordHelpKeywordui_login_tunnelCaptionTun
ImageIndex
TabVisible
DesignSizea  	TGroupBoxTunnelSessionGroupLeft Top WidthYHeight� AnchorsakLeftakTopakRight CaptionV�rd f�r att s�tta upp tunnelTabOrder
DesignSizeY�   TLabelLabel6LeftTopWidth6HeightCaption
&V�rdnamn:FocusControlTunnelHostNameEdit  TLabelLabel14Left� TopWidth<HeightAnchorsakTopakRight CaptionPo&rtnummer:FocusControlTunnelPortNumberEdit  TLabelLabel15LeftTopDWidth6HeightCaption&Anv�ndarnamn:FocusControlTunnelUserNameEdit  TLabelLabel16Left� TopDWidth1HeightCaption
&L�senord:FocusControlTunnelPasswordEdit  TLabelLabel18LeftTopvWidthHHeightCaptionFil med privat nyc&kelFocusControlTunnelPrivateKeyEdit  TEditTunnelHostNameEditLeftTop#Width� HeightAnchorsakLeftakTopakRight 	MaxLengthdTabOrder TextTunnelHostNameEditOnChange
DataChange  TEditTunnelUserNameEditLeftTopUWidth� Height	MaxLength2TabOrderTextTunnelUserNameEditOnChange
DataChange  TPasswordEditTunnelPasswordEditLeft� TopUWidth� HeightAnchorsakLeftakTopakRight 	MaxLength2TabOrderTextTunnelPasswordEditOnChange
DataChange  TUpDownEditTunnelPortNumberEditLeft� Top#WidthRHeight	AlignmenttaRightJustifyMaxValue��  MinValueValueAnchorsakTopakRight TabOrderOnChange
DataChange  TFilenameEditTunnelPrivateKeyEditLeftTop� WidthBHeightAcceptFiles	OnAfterDialogPrivateKeyEditAfterDialogFilter8PuTTY privata nycklar (*.ppk)|*.ppk|Alla filer (*.*)|*.*DialogOptions
ofReadOnlyofPathMustExistofFileMustExist DialogTitleV�lj fil med privat nyckelClickKey@AnchorsakLeftakTopakRight TabOrderTextTunnelPrivateKeyEditOnChange
DataChange   	TCheckBoxTunnelCheckLeftTopWidth3HeightCaptionAnslut med SSH-tunnelTabOrder OnClick
DataChange  	TGroupBoxTunnelOptionsGroupLeft Top� WidthYHeight/AnchorsakLeftakTopakRight CaptionAlternativ f�r tunnelTabOrder
DesignSizeY/  TLabelLabel21LeftTopWidthRHeightCaption&Lokal tunnelport:FocusControlTunnelLocalPortNumberEdit  	TComboBoxTunnelLocalPortNumberEditLeft� TopWidthRHeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeight	MaxLength2TabOrder TextTunnelLocalPortNumberEditOnChange
DataChangeItems.StringsV�lj automatiskt     	TTabSheetAdvancedSheetTagHintSSHHelpType	htKeywordHelpKeywordui_login_sshCaptionSSH
ImageIndex
TabVisible
DesignSizea  	TGroupBoxProtocolGroupLeft TopWidthYHeightWAnchorsakLeftakTopakRight CaptionAlternativ f�r protokollTabOrder 
DesignSizeYW  TLabelLabel7LeftTop*Width� HeightCaptionF�redragen SSH-version:FocusControlSshProt1onlyButton  TRadioButtonSshProt1ButtonLeftXTop;WidthAHeightCaption&1TabOrderOnClick
DataChange  TRadioButtonSshProt2ButtonLeft� Top;WidthAHeightCaption&2TabOrderOnClick
DataChange  	TCheckBoxCompressionCheckLeftTopWidthDHeightAnchorsakLeftakTopakRight CaptionAnv�nd &komprimeringTabOrder OnClick
DataChange  TRadioButtonSshProt1onlyButtonLeftTop;WidthAHeightCaption	End&ast 1Checked	TabOrderTabStop	OnClick
DataChange  TRadioButtonSshProt2onlyButtonLeft� Top;WidthAHeightCaption	&Endast 2TabOrderOnClick
DataChange   	TGroupBoxEncryptionGroupLeft TopdWidthYHeight� AnchorsakLeftakTopakRight CaptionKrypteringsinst�llningarTabOrder
DesignSizeY�   TLabelLabel8LeftTopWidth� HeightCaption#&Riktlinjer f�r krypteringschiffer:FocusControlCipherListBox  TListBoxCipherListBoxLeftTop$Width� Height[DragModedmAutomatic
ItemHeightTabOrder OnClick
DataChange
OnDragDropAlgListBoxDragDrop
OnDragOverAlgListBoxDragOverOnStartDragAlgListBoxStartDrag  	TCheckBoxSsh2LegacyDESCheckLeftTop� Width=HeightAnchorsakLeftakTopakRight Caption+Till�t arvsanv�nding av single-&DES i SSH-2TabOrder  TButtonCipherUpButtonLeft� Top$WidthFHeightCaption&UppTabOrderOnClickCipherButtonClick  TButtonCipherDownButtonLeft� TopDWidthFHeightCaption&NerTabOrderOnClickCipherButtonClick    	TTabSheetKexSheetTagHint
NyckelbyteHelpType	htKeywordHelpKeywordui_login_kexCaptionKEX
ImageIndex
TabVisible
DesignSizea  	TGroupBoxKexOptionsGroupLeft TopWidthYHeight� AnchorsakLeftakTopakRight Caption$Alternativ f�r nyckelbytesalgoritmenTabOrder  TLabelLabel28LeftTopWidthyHeightCaptionRi&ktlinjer f�r algoritmen:FocusControl
KexListBox  TListBox
KexListBoxLeftTop$Width� HeightYDragModedmAutomatic
ItemHeightTabOrder OnClick
DataChange
OnDragDropAlgListBoxDragDrop
OnDragOverAlgListBoxDragOverOnStartDragAlgListBoxStartDrag  TButtonKexUpButtonLeft� Top$WidthFHeightCaption&UppTabOrderOnClickKexButtonClick  TButtonKexDownButtonLeft� TopDWidthFHeightCaption&NerTabOrderOnClickKexButtonClick   	TGroupBoxKexReexchangeGroupLeft Top� WidthYHeightEAnchorsakLeftakTopakRight Caption'Alternativ f�r kontroll av nyckelutbyteTabOrder TLabelLabel31LeftTopWidth� HeightCaption>Max antal minuter innan nyckeluppdatering (0 ger ingen gr�ns):Color	clBtnFaceFocusControlRekeyTimeEditParentColor  TLabelLabel32LeftTop,Width� HeightCaption;Max antal data innan nyckeluppdatering (0 ger ingen gr�ns):Color	clBtnFaceFocusControlRekeyDataEditParentColor  TUpDownEditRekeyTimeEditLeft TopWidthIHeight	AlignmenttaRightJustifyMaxValue�	MaxLengthTabOrder OnChange
DataChange  TEditRekeyDataEditLeft Top'WidthIHeight	MaxLength
TabOrderOnChange
DataChange    	TTabSheet	AuthSheetTagHintAutentiseringHelpType	htKeywordHelpKeywordui_login_authenticationCaptionAuth
ImageIndex

TabVisible
DesignSizea  	TCheckBoxSshNoUserAuthCheckLeftTopWidth3HeightCaption-Kringg� autentisering helt och h�llet (SSH-2)TabOrder OnClick
DataChange  	TGroupBoxAuthenticationGroupLeft Top WidthYHeight� AnchorsakLeftakTopakRight CaptionAlternativ f�r autentiseringTabOrder
DesignSizeY�   	TCheckBoxTryAgentCheckLeftTopWidthEHeightAnchorsakLeftakTopakRight Caption)F�rs�k anv�nda autentisering med &PageantTabOrder OnClick
DataChange  	TCheckBoxAuthTISCheckLeftTop*WidthEHeightAnchorsakLeftakTopakRight Caption:F�rs�k anv�nda &TIS eller Kryptokort autentisering (SSH-1)TabOrderOnClick
DataChange  	TCheckBoxAuthKICheckLeftTopAWidthEHeightAnchorsakLeftakTopakRight Caption=F�rs�k anv�nda 'tagentbords&interaktiv' autentisering (SSH-2)TabOrderOnClick
DataChange  	TCheckBoxAuthKIPasswordCheckLeft TopXWidth1HeightAnchorsakLeftakTopakRight Caption'Svara med l�senord vid f�rsta &promptenTabOrderOnClick
DataChange  	TCheckBoxAuthGSSAPICheck2LeftTopoWidthEHeightCaption0F�rs�k anv�nda GSSAPI/SSPI autentisering (SSH-2)TabOrderOnClickAuthGSSAPICheck2Click   	TGroupBoxAuthenticationParamsGroupLeft Top� WidthYHeight0AnchorsakLeftakTopakRight CaptionParametrar autentiseringTabOrder
DesignSizeY0  	TCheckBoxAgentFwdCheckLeftTopWidthEHeightAnchorsakLeftakTopakRight CaptionTill�t agent-vidarebe&fordranTabOrder OnClick
DataChange    	TTabSheet	BugsSheetTagHintBuggarHelpType	htKeywordHelpKeywordui_login_bugsCaptionBugs
ImageIndex	
TabVisible
DesignSizea  	TGroupBoxBugsGroupBoxLeft TopWidthYHeight� AnchorsakLeftakTopakRight CaptionUppt�cka buggar i SSH-servrarTabOrder 
DesignSizeY�   TLabelBugIgnore1LabelLeftTopWidth� HeightCaption'Stannar vid &ignore-meddelanden i SSH-1FocusControlBugIgnore1Combo  TLabelBugPlainPW1LabelLeftTop,Width� HeightCaption'&V�grar all l�senordskamouflage i SSH1-FocusControlBugPlainPW1Combo  TLabelBugRSA1LabelLeftTopDWidth� HeightCaption&Stannar vid &RSA-autentisering i SSH-1FocusControlBugRSA1Combo  TLabelBugHMAC2LabelLeftTop\Width� HeightCaption&Ber�kningsfel av H&MAC-nycklar i SSH-2FocusControlBugHMAC2Combo  TLabelBugDeriveKey2LabelLeftToptWidth� HeightCaption,Ber�kningsf&el av krypteringsnycklar i SSH-2FocusControlBugDeriveKey2Combo  TLabelBugRSAPad2LabelLeftTop� Width� HeightCaption+Kr�ver &utfyllnad av RSA-signaturer i SSH-2FocusControlBugRSAPad2Combo  TLabelBugPKSessID2LabelLeftTop� Width� HeightCaption0Sessio&ns-id i SSH-2 PK autentisering missbrukasFocusControlBugPKSessID2Combo  TLabelBugRekey2LabelLeftTop� Width� HeightCaption$Hanterar SSH-2 nyc&kelutbyte d�ligt:FocusControlBugRekey2Combo  TLabelBugMaxPkt2LabelLeftTop� Width� HeightCaption*Ignorerar SSH-2 ma&ximum f�r paketstorlek:FocusControlBugMaxPkt2Combo  	TComboBoxBugIgnore1ComboLeftTopWidth=HeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrder OnChange
DataChange  	TComboBoxBugPlainPW1ComboLeftTop'Width=HeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrderOnChange
DataChange  	TComboBoxBugRSA1ComboLeftTop?Width=HeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrderOnChange
DataChange  	TComboBoxBugHMAC2ComboLeftTopWWidth=HeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrderOnChange
DataChange  	TComboBoxBugDeriveKey2ComboLeftTopoWidth=HeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrderOnChange
DataChange  	TComboBoxBugRSAPad2ComboLeftTop� Width=HeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrderOnChange
DataChange  	TComboBoxBugPKSessID2ComboLeftTop� Width=HeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrderOnChange
DataChange  	TComboBoxBugRekey2ComboLeftTop� Width=HeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrderOnChange
DataChange  	TComboBoxBugMaxPkt2ComboLeftTop� Width=HeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrderOnChange
DataChange    	TTabSheetGeneralSheetTagHintInst�llningarHelpType	htKeywordHelpKeywordui_login_preferencesCaptionInt
ImageIndex
TabVisible TLabelLabel13LeftTop� WidthhHeightCaption�vriga inst�llningar:  TButtonPreferencesButtonLeft� Top� WidthZHeightCaption&Inst�llningar...TabOrderOnClickPreferencesButtonClick  �TGeneralSettingsFrameGeneralSettingsFrameLeft TopWidthYHeight� TabOrder 
DesignSizeY�   �	TGroupBoxInterfaceGroupWidthY
DesignSizeY�   �TLabelCommanderDescriptionLabel2Width�   �TLabelExplorerDescriptionLabelWidth�       TPanel	LeftPanelLeft Top Width� Height(AlignalLeft
BevelOuterbvNoneTabOrder 
DesignSize� (  	TTreeViewNavigationTreeLeftTop	Width� HeightAnchorsakLeftakTopakRightakBottom HideSelectionHotTrack	IndentReadOnly	ShowButtonsShowRootTabOrder OnChangeNavigationTreeChangeOnCollapsingNavigationTreeCollapsing
Items.Data
�     !               ����       SessionX)               ����        Stored sessionsX!               ����        LoggingX%               ����       EnvironmentX%               ����        DirectoriesX%               ����        Recycle binX               ����        SFTPX               ����        SCPX           ��������        FTPX$               ����       ConnectionX               ����        ProxyX                ����        TunnelX               ����       SSHX&               ����        Kex exchangeX(               ����        AuthenticationX               ����        BugsX%               ����        PreferencesX  	TCheckBoxShowAdvancedLoginOptionsCheckLeftTopWidthxHeightAnchorsakLeftakRightakBottom Caption
&AvanceratTabOrderOnClick
DataChange    TActionList
ActionListOnUpdateActionListUpdateLeftTop TActionEditSessionActionCategorySessionsCaption	&Redigera	OnExecuteEditSessionActionExecute  TActionSaveSessionActionCategorySessionsCaption	&Spara...	OnExecuteSaveSessionActionExecute  TActionDeleteSessionActionCategorySessionsCaptionTa &bort...	OnExecuteDeleteSessionActionExecute  TActionImportSessionsActionCategorySessionsCaption&Importera...	OnExecuteImportSessionsActionExecute  TActionLoginActionCategorySessionCaptionLogga in  TActionAboutActionCategoryOtherCaption&Om...	OnExecuteAboutActionExecute  TActionCleanUpActionCategoryOtherCaption&Rensa applikationsdata...	OnExecuteCleanUpActionExecute  TActionNewSessionActionCategorySessionsCaption&Ny	OnExecuteNewSessionActionExecute  TActionSetDefaultSessionActionCategorySessionsCaptionS�&tt standard	OnExecuteSetDefaultSessionActionExecute  TActionDesktopIconActionCategorySessionsCaptionSkrivbords&ikon	OnExecuteDesktopIconActionExecute  TActionSendToHookActionCategorySessionsCaption!Utforskarens 'Skicka till'-genv�g	OnExecuteSendToHookActionExecute  TActionCheckForUpdatesActionTagCategoryOtherCaptionS�k efter &uppdateringar
ImageIndex?	OnExecuteCheckForUpdatesActionExecute  TActionRenameSessionActionCategorySessionsCaption	Byt &namn	OnExecuteRenameSessionActionExecute  TActionShellIconSessionActionCategorySessionsCaption	Skal&ikon	OnExecuteShellIconSessionActionExecute  TActionNewSessionFolderActionCategorySessionsCaptionN&y mapp...	OnExecuteNewSessionFolderActionExecute   
TPopupMenuToolsPopupMenuLeft0Top 	TMenuItemImport1ActionImportSessionsAction  	TMenuItemCleanup1ActionCleanUpAction  	TMenuItemCheckForUpdates1ActionCheckForUpdatesAction   
TPopupMenuIconsPopupMenuLeftPTop 	TMenuItemDesktopicon1ActionDesktopIconAction  	TMenuItemExplorersSendtoshortcut1ActionSendToHookAction   
TPopupMenuColorPopupMenuImagesColorImageListLeftpTop 	TMenuItemColorDefaultItemCaption	&StandardOnClickColorDefaultItemClick  	TMenuItemPickColorItemCaption&V�lj f�rg...
ImageIndex OnClickPickColorItemClick   
TImageListColorImageListBkColorclRedAllocByLeftTop!Bitmap
&  IL     �   ���������BM6       6   (   @                                  �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                 BM>       >   (   @            �                       ��� ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��                              
TImageListSessionImageListLeft0Top!Bitmap
&2  IL 	    �������������BM6       6   (   @   0           0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              !! !! !! !! !! !! !! !! !! !! !! !!                                                                                                                                                                                                              cc  cc  cc  cc  cc  cc  cc  cc  cc  cc  cc !! !!          cc ���  ��  ��  ��  ��  ��  ��  ��  ��  �� c��  ��                                                                                                                                                  cc ���  ��  ��  ��  ��  ��  ��  ��  ��  cc !! !!          cc ���  ��  ��  ��  ��  ��  ��  ��  ��  ��  �� c��                                                                                                                                              cc ���  ��  ��  ��  ��  ��  ��  ��  �� c�� !!  cc !!          cc ��� ���  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��                                                                                                                                              cc ��� ���  ��  ��  ��  ��  ��  ��  ��  �� !!  cc !!          cc ���  �� ���  ��  ��  ��  ��  ��  ��  ��  ��  ��                                                                                                                                          cc ��� ���  �� ���  ��  ��  ��  ��  ��  �� !!  ��  �� !!          cc ��� ���  �� ���  ��  ��  ��  ��  ��  ��  ��  ��                                                                                                                                          cc ���  �� ���  �� ���  ��  ��  ��  ��  �� !!  ��  �� !!          cc ���  �� ���  �� ���  �� ���  ��  ��  ��  ��  ��                                                                                                                                          cc  cc  cc  cc  cc  cc  cc  cc  cc  cc  cc  ��  ��  �� !!          cc ��� ���  �� ���  �� ���  �� ���  ��  ��  ��  ��                                                                                                                                              cc ���  �� ���  ��  ��  ��  ��  ��  ��  ��  ��  �� !!          cc ���  �� ���  �� ���  �� ���  �� ���  ��  ��  ��                                                                                                                                              cc ��� ���  �� ���  ��  ��  ��  �� ��� ��� ��� ��� !!          cc ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                                                                              cc ���  �� ���  �� ���  �� ���  cc  cc  cc  cc  cc              cc  cc  cc  cc  cc  cc  cc  cc  cc  cc  cc  cc  cc                                                                                                                                                  cc ��� ��� ��� ��� ���  cc                                      cc ��� ��� ��� ���  ��                                                                                                                                                                              cc  cc  cc  cc  cc                                              cc  cc  cc  cc  cc                                                                                                                                                                                                                                                                                                 BM>       >   (   @   0         �                      ���                                                                                                                                                                                                                                                                 �������������������������������������������������� ����� ����� �����������������������������������������                           TPF0TNonVisualDataModuleNonVisualDataModuleOldCreateOrderLeftTop� Height�Widthp TActionList
LogActionsImagesGlyphsModule.LogImages	OnExecuteLogActionsExecuteOnUpdateLogActionsUpdateLeft Toph TActionLogClearActionCategoryLogMemoCaption&RensaHint
Rensa logg
ImageIndexShortCut.@  TActionLogSelectAllActionCategoryLogMemoCaptionM&arkera alltHintMarkera allt
ImageIndexShortCutA@  TActionLogCopyActionCategoryLogMemoCaption&KopieraHintKopiera till urklipp
ImageIndexShortCutC@  TActionLogCloseActionCategoryLogFormCaptionSt&�ngHintSt�ng loggf�nster
ImageIndex ShortCuts�    TActionLogPreferencesActionCategoryLogFormCaptionLogPreferencesActionHintKonfigurera loggning
ImageIndex   TTBXPopupMenuLogMemoPopupImagesGlyphsModule.LogImagesLeft Top�  TTBXItemClear1ActionLogClearAction  TTBXItemClose1ActionLogCopyAction  TTBXItem
Selectall1ActionLogSelectAllAction   TTBXPopupMenuRemoteFilePopupImagesGlyphsModule.ExplorerImagesLeft�TopP TTBXItem	TBXItem23ActionAddEditLinkContextAction  TTBXItemCurrentOpenMenuItemActionCurrentOpenAction  TTBXItemCurrentEditMenuItemActionCurrentEditFocusedAction  TTBXItemCurrentCopyMenuItemActionCurrentCopyFocusedAction  TTBXItem
Duplicate3ActionRemoteCopyToAction  TTBXItemMoveto1ActionCurrentMoveFocusedAction  TTBXItemMoveto6ActionRemoteMoveToFocusedAction  TTBXItemDelete1ActionCurrentDeleteFocusedAction  TTBXItemRename1ActionCurrentRenameAction  TTBXSeparatorItemN45  TTBXSubmenuItemRemoteDirViewCustomCommandsMenuActionCustomCommandsAction TTBXItem    TTBXSubmenuItem
FileNames3Caption&FilnamnHelpKeyword	filenamesHint'Operationer med namn p� vald(a) fil(er) TTBXItemInserttoCommandLine2ActionFileListToCommandLineAction  TTBXItemCopytoClipboard3ActionFileListToClipboardAction  TTBXItemCopytoClipboardIncludePaths3ActionFullFileListToClipboardAction  TTBXItemCopyURLtoClipboard3ActionUrlToClipboardAction   TTBXSeparatorItemN1  TTBXItemProperties1ActionCurrentPropertiesFocusedAction   TActionListExplorerActionsImagesGlyphsModule.ExplorerImages	OnExecuteExplorerActionsExecuteOnUpdateExplorerActionsUpdateLeft�Top TActionBestFitColumnActionTagCategoryColumnsCaption&B�sta passningHint4B�sta passning|Anpassa kolumnbredden till inneh�llet  TActionGoToTreeActionTagCategoryViewCaptionG� till tr�dHelpKeywordui_file_panel#directory_treeHintG� till tr�d
ImageIndexLShortCutT�    TActionLocalTreeActionTagCategoryViewCaption&Tr�dHelpKeywordui_file_panel#directory_treeHintD�lj/visa katalogtr�d
ImageIndexLShortCutT�    TActionRemoteTreeActionTagCategoryViewCaption&Tr�dHelpKeywordui_file_panel#directory_treeHintD�lj/visa katalogtr�d
ImageIndexLShortCutT�    TActionQueueItemQueryActionTagCategoryQueueCaptionVi&sa fr�gaHelpKeywordui_queue#managing_the_queueHint$Visa avvaktande fr�ga p� vald k�post
ImageIndexC  TActionQueueItemErrorActionTagCategoryQueueCaption	Vi&sa felHelpKeywordui_queue#managing_the_queueHint,Visa avvaktande felmeddelande p� vald k�post
ImageIndexD  TActionQueueItemPromptActionTagCategoryQueueCaptionVi&sa promptHelpKeywordui_queue#managing_the_queueHint%Visa avvaktande prompt p� vald k�post
ImageIndexE  TActionGoToCommandLineActionTagCategoryViewCaptionG� till komma&ndoradHelpKeywordui_commander#command_lineHintG� till kommandoradShortCutN`  TActionQueueItemDeleteActionTagCategoryQueueCaption&AvbrytHelpKeywordui_queue#managing_the_queueHintTa bort vald k�post
ImageIndexG  TActionQueueItemExecuteActionTagCategoryQueueCaption	&Utf�r nuHelpKeywordui_queue#managing_the_queueHintAUtf�r vald k�post omedelbart genom att ge den en extra anslutning
ImageIndexF  TActionSelectOneActionTagCategory	SelectionCaption&Markera/avmarkeraHelpKeywordui_file_panel#selecting_filesHint"Markera|Markera/avmarkera vald fil  TActionCurrentRenameActionTagCategory5Toolbar Operation (selected + rename + mkdir + close)Caption	&Byt namnHelpKeywordtask_renameHintByt namn|Byt namn p� vald fil
ImageIndex  TActionLocalSortAscendingActionTag	CategorySortCaption	Stig&andeHelpKeywordui_file_panel#sorting_filesHintSStigande/fallande|V�xla mellan stigande och fallande sortering i den lokala panelen
ImageIndex%  TActionCurrentEditActionTagCategory5Toolbar Operation (selected + rename + mkdir + close)Caption	&RedigeraHelpKeyword	task_editHintRedigera|Redigera markerad fil
ImageIndex9  TActionHideColumnActionTagCategoryColumnsCaption&D�lj kolumnHelpKeywordui_file_panel#selecting_columnsHintD�lj kolumn|D�lj vald kolumn  TActionLocalBackActionTag	CategoryLocal DirectoryCaption	Till&bakaHelpKeywordtask_navigate#special_commands
ImageIndexShortCut%�    TActionCurrentCopyActionTagCategory5Toolbar Operation (selected + rename + mkdir + close)CaptionK&opiera...HelpKeywordtask_downloadHintKopiera|Kopiera markerade filer
ImageIndex   TActionCurrentMoveActionTagCategory5Toolbar Operation (selected + rename + mkdir + close)Caption
&Flytta...HelpKeywordtask_downloadHintFlytta|Flytta markerade filer
ImageIndex  TActionCurrentCycleStyleActionTagCategoryStyleCaptionVisaHelpKeywordui_file_panel#view_styleHint7Visa|V�xla mellan att visa olika stilar f�r katalogvyer
ImageIndex  TActionCurrentIconActionTagCategoryStyleCaptionSt&ora ikonerHelpKeywordui_file_panel#view_styleHintStora ikoner|Visa stora ikoner
ImageIndex  TActionCurrentSmallIconActionTagCategoryStyleCaption&Sm� ikonerHelpKeywordui_file_panel#view_styleHintSm� ikoner|Visa sm� ikoner
ImageIndex	  TActionCurrentListActionTagCategoryStyleCaptionLis&taHelpKeywordui_file_panel#view_styleHintLista|Visa lista
ImageIndex
  TActionCurrentReportActionTagCategoryStyleCaption&Detaljerad listaHelpKeywordui_file_panel#view_styleHint&Detaljerad lista|Visa detaljerad lista
ImageIndex  TActionCurrentCopyFocusedActionTagCategoryFocused OperationCaptionK&opiera...HelpKeywordtask_downloadHint2Kopiera|Kopiera markerade filer till lokal katalog
ImageIndex   TActionRemoteMoveToActionTagCategorySelected OperationCaption&Flytta till...HelpKeyword'task_move_duplicate#moving_remote_filesHint/Flytta|Flytta markerade filer till fj�rrkatalog  TActionCurrentMoveFocusedActionTagCategoryFocused OperationCaption
&Flytta...HelpKeywordtask_downloadHint0Flytta|Flytta markerade filer till lokal katalog
ImageIndex  TActionCurrentDeleteFocusedActionTagCategoryFocused OperationCaption&Ta bortHelpKeywordtask_deleteHintTa bort|Ta bort markerade filer
ImageIndex  TActionCurrentPropertiesFocusedActionTagCategoryFocused OperationCaption&EgenskaperHelpKeywordtask_propertiesHint4Egenskaper|Visa/�ndra egenskaper f�r markerade filer
ImageIndex  TActionCurrentCreateDirActionTagCategory5Toolbar Operation (selected + rename + mkdir + close)CaptionS&kapa katalog...HelpKeywordtask_create_directoryHintSkapa katalog|Skapa ny katalog
ImageIndex  TActionCurrentDeleteActionTagCategory5Toolbar Operation (selected + rename + mkdir + close)Caption&Ta bortHelpKeywordtask_deleteHintTa bort|Ta bort markerade filer
ImageIndex  TActionCurrentPropertiesActionTagCategory5Toolbar Operation (selected + rename + mkdir + close)Caption&EgenskaperHelpKeywordtask_propertiesHint4Egenskaper|Visa/�ndra egenskaper f�r markerade filer
ImageIndex  TActionRemoteBackActionTagCategoryRemote DirectoryCaption	Till&bakaHelpKeywordtask_navigate#special_commands
ImageIndexShortCut%�    TActionRemoteForwardActionTagCategoryRemote DirectoryCaption&Fram�tHelpKeywordtask_navigate#special_commands
ImageIndexShortCut'�    TActionCommandLinePanelActionTagCategoryViewCaptionKomma&ndoradHelpKeywordui_commander#command_lineHintD�lj/visa kommandoradShortCutN`  TActionRemoteParentDirActionTagCategoryRemote DirectoryCaption&�verliggande katalogHelpKeywordtask_navigate#special_commandsHint!Huvudkatalog|G� till huvudkatalog
ImageIndex  TActionRemoteRootDirActionTagCategoryRemote DirectoryCaption&RotkatalogHelpKeywordtask_navigate#special_commandsHintRotkatalog|G� till rotkatalog
ImageIndexShortCut�@  TActionRemoteHomeDirActionTagCategoryRemote DirectoryCaption&HemkatalogHelpKeywordtask_navigate#special_commandsHintHemkatalog|G� till hemkatalog
ImageIndex  TActionRemoteRefreshActionTagCategoryRemote DirectoryCaption
&UppdateraHint#Uppdatera|Uppdatera kataloginneh�ll
ImageIndex  TActionAboutActionTagCategoryHelpCaption&Om...HelpKeywordui_aboutHintOm|Visa programinformation
ImageIndex  TActionStatusBarActionTagCategoryViewCaption&Statusf�ltHintVisa/d�lj statusf�ltet  TActionExplorerAddressBandActionTagCategoryViewCaption&AdressHelpKeywordui_toolbarsHintVisa/d�lj adressf�ltet  TActionExplorerMenuBandActionTagCategoryViewCaption&MenyHelpKeywordui_toolbarsHintVisa/d�lj meny  TActionExplorerToolbarBandActionTagCategoryViewCaption&StandardknapparHelpKeywordui_toolbarsHint Visa/d�lj standardverktygsf�ltet  TActionRemoteOpenDirActionTagCategoryRemote DirectoryCaption&�ppna katalog/bokm�rkeHelpKeyword$task_navigate#entering_path_manuallyHint?�ppna katalog/bokm�rke|�ppna vald katalog eller sparat bokm�rke
ImageIndex  TActionSelectActionTagCategory	SelectionCaption&Markera filerHelpKeyword	ui_selectHint)Markera|Markera filer beroende p� filmask
ImageIndex  TActionUnselectActionTagCategory	SelectionCaptionA&vmarkera filerHelpKeyword	ui_selectHint-Avmarkera|Avmarkera filer beroende p� filmask
ImageIndex  TActionSelectAllActionTagCategory	SelectionCaptionM&arkera allaHelpKeywordui_file_panel#selecting_filesHintMarkera alla
ImageIndex  TActionInvertSelectionActionTagCategory	SelectionCaption&Inverterad markeringHelpKeywordui_file_panel#selecting_filesHintInverterad markering
ImageIndex  TActionExplorerSelectionBandActionTagCategoryViewCaption&MarkeringsknapparHelpKeywordui_toolbarsHint&D�lj/visa verktygsf�ltet f�r markering  TActionClearSelectionActionTagCategory	SelectionCaption&Rensa markeringHelpKeywordui_file_panel#selecting_filesHintRensa markering
ImageIndex  TActionExplorerSessionBandActionTagCategoryViewCaptionSessio&nsknapparHelpKeywordui_toolbarsHint&D�lj/visa verktygsf�ltet f�r sessioner  TActionExplorerPreferencesBandActionTagCategoryViewCaptionInst�llningsknapparHelpKeywordui_toolbarsHint*Visa/d�lj verktygsf�ltet f�r inst�llningar  TActionExplorerSortBandActionTagCategoryViewCaptionSo&rteringsknapparHelpKeywordui_toolbarsHint&Visa/d�lj verktygsf�ltet f�r sortering  TActionExplorerUpdatesBandActionTagCategoryViewCaption&UppdateringknappHelpKeywordui_toolbarsHint)D�lj/visa verktykgsf�lt f�r uppdateringar  TActionExplorerTransferBandActionTagCategoryViewCaption&�verf�r inst�llningarHelpKeywordui_toolbarsHint3D�lj/visa verktygsf�lt f�r �verf�ringsinst�llningar  TAction ExplorerCustomCommandsBandActionTagCategoryViewCaptionEgna ko&mmandoknapparHelpKeywordui_toolbarsHint)D�lj/visa verktygsf�lt f�r egna kommandon  TActionViewLogActionTagCategoryViewCaptionLo&ggf�nsterHelpKeywordui_logHintVisa/d�lj loggf�nster
ImageIndex  TActionNewSessionActionTagCategorySessionCaption&Ny session...HelpKeyword.task_connections#opening_additional_connectionHintRNy session|�ppna ny session (H�ll nere SHIFT f�r att �ppna den i ett nytt f�nster)
ImageIndexShortCutN@SecondaryShortCuts.StringsCtrl+Shift+N   TActionCloseSessionActionTagCategorySessionCaption&Koppla ifr�nHint%St�ng session|Avsluta aktuell session
ImageIndexShortCutD`  TActionSavedSessionsActionTagCategorySessionCaptionS&parade sessionerHelpKeyword.task_connections#opening_additional_connectionHint�ppna sparad session
ImageIndex  TActionPreferencesActionTagCategoryViewCaption&Inst�llningar...HelpKeywordui_preferencesHint.Inst�llningar|Visa/�ndra anv�ndarinst�llningar
ImageIndexShortCutP�    TActionRemoteChangePathActionTagCategoryRemote DirectoryCaption&Byt katalogHelpKeywordtask_navigateHint.Till�ter att annan katalog v�lj i fj�rrpanelen
ImageIndexShortCutq�    TActionLocalForwardActionTag	CategoryLocal DirectoryCaption&Fram�tHelpKeywordtask_navigate#special_commands
ImageIndexShortCut'�    TActionLocalParentDirActionTagCategoryLocal DirectoryCaption&HuvudkatalogHelpKeywordtask_navigate#special_commandsHint!Huvudkatalog|G� till huvudkatalog
ImageIndex  TActionLocalRootDirActionTagCategoryLocal DirectoryCaption&RotkatalogHelpKeywordtask_navigate#special_commandsHintRotkatalog|G� till rotkatalogen
ImageIndexShortCut�@  TActionLocalHomeDirActionTag	CategoryLocal DirectoryCaption&HemkatalogHelpKeywordtask_navigate#special_commandsHintHemkatalog|G� till hemkatalogen
ImageIndex  TActionLocalRefreshActionTag	CategoryLocal DirectoryCaption
&UppdateraHint#Uppdatera|Uppdatera kataloginneh�ll
ImageIndex  TActionLocalOpenDirActionTag	CategoryLocal DirectoryCaption&�ppna katalog/bokm�rke...HelpKeyword$task_navigate#entering_path_manuallyHint?�ppna katalog/bokm�rke|�ppna vald katalog eller sparat bokm�rke
ImageIndex  TActionLocalChangePathActionTagCategoryLocal DirectoryCaption
&Byt enhetHelpKeywordtask_navigateHint.Till�ter att annan enhet v�ljs f�r lokal panel
ImageIndexShortCutp�    TActionToolBarActionTagCategoryViewCaptionKommandoverktygsf�ltHelpKeywordui_toolbarsHint$D�lj/visa verktygsf�lt f�r kommandon  TActionCommanderMenuBandActionTagCategoryViewCaption&MenyHelpKeywordui_toolbarsHintD�lj/visa meny  TActionCommanderSessionBandActionTagCategoryViewCaptionSessio&nsknapparHelpKeywordui_toolbarsHint&D�lj/visa verktygsf�ltet f�r sessioner  TActionCommanderPreferencesBandActionTagCategoryViewCaptionInst�llningsknapparHelpKeywordui_toolbarsHint*D�lj/visa verktygsf�ltet f�r inst�llningar  TActionCommanderSelectionBandActionTagCategoryViewCaption&MarkeringsknapparHelpKeywordui_toolbarsHint&D�lj/visa verktygsf�ltet f�r markering  TActionCommanderToolbarBandActionTagCategoryViewCaption&StandardknapparHelpKeywordui_toolbarsHint D�lj/visa standardverktygsf�ltet  TActionCommanderSortBandActionTagCategoryViewCaptionS&orteringsknapparHelpKeywordui_toolbarsHint&D�lj/visa verktygsf�ltet f�r sortering  TActionCommanderUpdatesBandActionTagCategoryViewCaption&UppdateringsknappHelpKeywordui_toolbarsHint&D�lj/visa verktygsf�lt f�r uppdatering  TActionCommanderTransferBandActionTagCategoryViewCaption�verf�ringsinst�llningarHelpKeywordui_toolbarsHint3D�lj/visa verktygsf�lt f�r �verf�ringsinst�llningar  TActionCommanderCommandsBandActionTagCategoryViewCaption&KommandoknapparHelpKeywordui_toolbarsHint&Visa/d�lj verktygsf�ltet f�r kommandon  TAction!CommanderUploadDownloadBandActionTagCategoryViewCaptionUp&p/nerladdningsknapparHelpKeywordui_toolbarsHint*D�lj/visa verktygsf�lt f�r ner/uppladdning  TAction!CommanderCustomCommandsBandActionTagCategoryViewCaptionEgna ko&mmandoknapparHelpKeywordui_toolbarsHint)D�lj/visa verktygsf�lt f�r egna kommandon  TActionCommanderLocalHistoryBandActionTagCategoryViewCaption&HistorikknapparHelpKeywordui_toolbarsHint+D�lj/visa verktygsf�ltet f�r lokal historik  TAction"CommanderLocalNavigationBandActionTagCategoryViewCaption&NavigeringsknapparHelpKeywordui_toolbarsHint-D�lj/visa verktygsf�ltet f�r lokal navigering  TAction CommanderRemoteHistoryBandActionTagCategoryViewCaption&HistorikknapparHelpKeywordui_toolbarsHint&D�lj/visa verktygsf�ltet fj�rrhistorik  TAction#CommanderRemoteNavigationBandActionTagCategoryViewCaption&NavigeringsknapparHelpKeywordui_toolbarsHint,D�lj/visa verktygsf�ltet f�r fj�rrnavigering  TActionLocalStatusBarActionTagCategoryViewCaptionStatusf&�ltHint(D�lj/visa den lokala panelens statusf�lt  TActionRemoteStatusBarActionTagCategoryViewCaptionStatusf&�ltHint"D�lj/visa fj�rrpanelens statusf�lt  TActionLocalSortByNameActionTag	CategorySortCaptionEfter &namnHelpKeywordui_file_panel#sorting_filesHint8Sortera efter namn|Sortera den lokala panelen efter namn
ImageIndexShortCutr@  TActionLocalSortByExtActionTag	CategorySortCaptionEfter &fil�ndelseHelpKeywordui_file_panel#sorting_filesHintDSortera efter fil�ndelse|Sortera den lokala panelen efter fil�ndelse
ImageIndex ShortCuts@  TActionLocalSortBySizeActionTag	CategorySortCaptionEfter &storlekHelpKeywordui_file_panel#sorting_filesHintASortera efter storlek|Sortera den lokala panelen efter filstorlek
ImageIndex#ShortCutu@  TActionLocalSortByAttrActionTag	CategorySortCaptionEfter &attributHelpKeywordui_file_panel#sorting_filesHint@Sortera efter attribut|Sortera den lokala panelen efter attribut
ImageIndex$ShortCutv@  TActionLocalSortByTypeActionTag	CategorySortCaptionEfter fil&typHelpKeywordui_file_panel#sorting_filesHint<Sortera efter filtyp|Sortera den lokala panelen efter filtyp
ImageIndex"  TActionLocalSortByChangedActionTag	CategorySortCaptionEfter senast &�ndradHelpKeywordui_file_panel#sorting_filesHintKSortera efter senast &�ndrad|Sortera den lokala panelen efter senast �ndrad
ImageIndex!ShortCutt@  TActionRemoteSortAscendingActionTagCategorySortCaption	Stig&andeHelpKeywordui_file_panel#sorting_filesHintUStigande/fallande|V�xla sortering mellan stigande och fallande ordning i fj�rrpanelen
ImageIndex%  TActionRemoteSortByNameActionTagCategorySortCaptionEfter &namnHelpKeywordui_file_panel#sorting_filesHint2Sortera efter namn|Sortera fj�rrpanelen efter namn
ImageIndexShortCutr@  TActionRemoteSortByExtActionTagCategorySortCaptionEfter &fil�ndelseHelpKeywordui_file_panel#sorting_filesHint>Sortera efter fil�ndelse|Sortera fj�rrpanelen efter fil�ndelse
ImageIndex ShortCuts@  TActionRemoteSortBySizeActionTagCategorySortCaptionEfter &storlekHelpKeywordui_file_panel#sorting_filesHint;Sortera efter storlek|Sortera fj�rrpanelen efter filstorlek
ImageIndex#ShortCutu@  TActionRemoteSortByRightsActionTagCategorySortCaptionEfter &filr�ttigheterHelpKeywordui_file_panel#sorting_filesHintFSortera efter filr�ttigheter|Sortera fj�rrpanelen efter filr�ttigheter
ImageIndex$ShortCutv@  TActionRemoteSortByChangedActionTagCategorySortCaptionEfter senast &�ndradHelpKeywordui_file_panel#sorting_filesHintESortera efter senast &�ndrad|Sortera fj�rrpanelen efter senast �ndrad
ImageIndex!ShortCutt@  TActionRemoteSortByOwnerActionTagCategorySortCaptionEfter �&gareHelpKeywordui_file_panel#sorting_filesHint7Sortera efter �gare|Sortera fj�rrpanelen efter fil�gare
ImageIndex&ShortCutw@  TActionRemoteSortByGroupActionTagCategorySortCaptionEfter &gruppHelpKeywordui_file_panel#sorting_filesHint7Sortera efter grupp|Sortera fj�rrpanelen efter filgrupp
ImageIndex'ShortCutx@  TActionRemoteSortByTypeActionTagCategorySortCaptionEfter fil&typHelpKeywordui_file_panel#sorting_filesHint6Sortera efter filtyp|Sortera fj�rrkatalog efter filtyp
ImageIndex"  TActionCurrentSortAscendingActionTagCategorySortCaption	Stig&andeHelpKeywordui_file_panel#sorting_filesHintVStigande/fallande|V�xla sortering mellan stigande och fallande ordning i aktuell panel
ImageIndex%  TActionCurrentSortByNameActionTagCategorySortCaptionEfter &namnHelpKeywordui_file_panel#sorting_filesHint3Sortera efter namn|Sortera aktuell panel efter namn
ImageIndexShortCutr@  TActionCurrentSortByExtActionTagCategorySortCaptionEfter &fil�ndelseHelpKeywordui_file_panel#sorting_filesHint?Sortera efter fil�ndelse|Sortera aktuell panel efter fil�ndelse
ImageIndex ShortCuts@  TActionCurrentSortBySizeActionTagCategorySortCaptionEfter &storlekHelpKeywordui_file_panel#sorting_filesHint<Sortera efter storlek|Sortera aktuell panel efter filstorlek
ImageIndex#ShortCutu@  TActionCurrentSortByTypeActionTagCategorySortCaptionEfter fil&typHelpKeywordui_file_panel#sorting_filesHintLSortera efter filtyp|Sortera aktuell panel efter filtyp (endast lokal panel)
ImageIndex"  TActionCurrentSortByRightsActionTagCategorySortCaptionEfter &attributHelpKeywordui_file_panel#sorting_filesHintJSortera efter attribut|Sortera aktuell panel efter attribut/filr�ttigheter
ImageIndex$ShortCutv@  TActionCurrentSortByChangedActionTagCategorySortCaptionEfter senast &�ndradHelpKeywordui_file_panel#sorting_filesHintFSortera efter senast &�ndrad|Sortera aktuell panel efter senast �ndrad
ImageIndex!ShortCutt@  TActionCurrentSortByOwnerActionTagCategorySortCaptionEfter �&gareHelpKeywordui_file_panel#sorting_filesHintLSortera efter �gare|Sortera aktuell panel efter fil�gare (endast fj�rrpanel)
ImageIndex&ShortCutw@  TActionCurrentSortByGroupActionTagCategorySortCaptionEfter &gruppHelpKeywordui_file_panel#sorting_filesHintKSortera efter grupp|Sortera fj�rrpanelen efter filgrupp (endast fj�rrpanel)
ImageIndex'ShortCutx@  TActionSortColumnAscendingActionTagCategorySortCaptionSortera stig&andeHelpKeywordui_file_panel#sorting_filesHint(Sortera filer stigande efter vald kolumn
ImageIndex)  TActionSortColumnDescendingActionTagCategorySortCaptionSortera fallan&deHelpKeywordui_file_panel#sorting_filesHint(Sortera filer fallande efter vald kolumn
ImageIndex(  TActionHomepageActionTagCategoryHelpCaptionProdukt&hemsidaHint6�ppnar webbl�saren och g�r till applikationens hemsida
ImageIndex*  TActionHistoryPageActionTagCategoryHelpCaption&VersionshistorikHintL�ppnar webbl�saren och g�r till webbsida med applikationens versionshistorik  TActionSaveCurrentSessionActionTagCategorySessionCaption&Spara session...HelpKeyword&task_connections#saving_opened_sessionHint#Spara session|Spara aktuell session
ImageIndex+  TActionShowHideRemoteNameColumnActionTagCategoryColumnsCaption&NamnHelpKeywordui_file_panel#selecting_columnsHint2Visa/d�lj namn|Visa/d�lj namnkolumn i fj�rrpanelen
ImageIndex,  TActionShowHideRemoteExtColumnActionTagCategoryColumnsCaption&Fil�ndelseHelpKeywordui_file_panel#selecting_columnsHint>Visa/d�lj fil�ndelse|Visa/d�lj fil�ndelsekolumn i fj�rrpanelen
ImageIndex-  TActionShowHideRemoteSizeColumnActionTagCategoryColumnsCaption&StorlekHelpKeywordui_file_panel#selecting_columnsHint<Visa/d�lj storlek|Visa/d�lj filstorlekskolumn i fj�rrpanelen
ImageIndex/  TAction!ShowHideRemoteChangedColumnActionTagCategoryColumnsCaptionSe&nast �ndradHelpKeywordui_file_panel#selecting_columnsHintEVisa/d�lj senast �ndrad|Visa/d�lj senast �ndrad-kolumn i fj�rrpanelen
ImageIndex0  TAction ShowHideRemoteRightsColumnActionTagCategoryColumnsCaptionFil&r�ttigheterHelpKeywordui_file_panel#selecting_columnsHintEVisa/d�lj filr�ttigheter|Visa/d�lj filr�ttighetskolumn i fj�rrpanelen
ImageIndex1  TActionShowHideRemoteOwnerColumnActionTagCategoryColumnsCaption&�gareHelpKeywordui_file_panel#selecting_columnsHint3Visa/d�lj �gare|Visa/d�lj �garkolumn i fj�rrpanelen
ImageIndex2  TActionShowHideRemoteGroupColumnActionTagCategoryColumnsCaption&GruppHelpKeywordui_file_panel#selecting_columnsHint4Visa/d�lj grupp|Visa/d�lj gruppkolumn i fj�rrpanelen
ImageIndex3  TAction$ShowHideRemoteLinkTargetColumnActionTagCategoryColumnsCaption&L�nkm�lHelpKeywordui_file_panel#selecting_columnsHint9Visa/d�lj l�nkm�l|Visa/d�lj l�nkm�lskolumn i fj�rrpanelen
ImageIndexR  TActionShowHideRemoteTypeColumnActionTagCategoryColumnsCaptionFil&typHelpKeywordui_file_panel#selecting_columnsHint7Visa/d�lj filtyp|Visa/d�lj filtypskolumn i fj�rrpanelen
ImageIndex.  TActionShowHideLocalNameColumnActionTagCategoryColumnsCaption&NamnHelpKeywordui_file_panel#selecting_columnsHint8Visa/d�lj namn|Visa/d�lj namnkolumn i den lokala panelen
ImageIndex,  TActionShowHideLocalExtColumnActionTagCategoryColumnsCaption&Fil�ndelseHelpKeywordui_file_panel#selecting_columnsHintDVisa/d�lj fil�ndelse|Visa/d�lj fil�ndelsekolumn i den lokala panelen
ImageIndex-  TActionShowHideLocalTypeColumnActionTagCategoryColumnsCaptionFil&typHelpKeywordui_file_panel#selecting_columnsHint=Visa/d�lj filtyp|Visa/d�lj filtypskolumn i den lokala panelen
ImageIndex.  TActionShowHideLocalSizeColumnActionTagCategoryColumnsCaption&StorlekHelpKeywordui_file_panel#selecting_columnsHintBVisa/d�lj storlek|Visa/d�lj filstorlekskolumn i den lokala panelen
ImageIndex/  TAction ShowHideLocalChangedColumnActionTagCategoryColumnsCaptionSenast &�ndradHelpKeywordui_file_panel#selecting_columnsHintKVisa/d�lj senast �ndrad|Visa/d�lj senast �ndrad-kolumn i den lokala panelen
ImageIndex0  TActionShowHideLocalAttrColumnActionTagCategoryColumnsCaption	&AttributHelpKeywordui_file_panel#selecting_columnsHint@Visa/d�lj attribut|Visa/d�lj attributkolumn i den lokala panelen
ImageIndex1  TActionCompareDirectoriesActionTagCategoryCommandCaption&J�mf�r katalogerHelpKeywordtask_compare_directoriesHintEJ�mf�r kataloger|Markerar skillnader mellan lokal- och fj�rrkatalogen
ImageIndex4ShortCutq   TActionSynchronizeActionTagCategoryCommandCaption&H�ll fj�rrkatalogen uppdateradHelpKeywordtask_keep_up_to_dateHint=H�ll fj�rrkatalogen uppdaterad|H�ll fj�rrkatalogen uppdaterad
ImageIndex5ShortCutU@  TActionForumPageActionTagCategoryHelpCaption&SupportforumHint:�ppnar webbl�saren och g� till webbsida med supportforumet  TActionLocalAddBookmarkActionTag	CategoryLocal DirectoryCaption&L�gg till bokm�rkenHelpKeywordtask_navigate#bookmarksHint@L�gg till bokm�rken|L�gg till aktuell lokal katalog som bokm�rke
ImageIndex6ShortCutB@  TActionRemoteAddBookmarkActionTagCategoryRemote DirectoryCaption&L�gg till bokm�rkenHelpKeywordtask_navigate#bookmarksHint?L�gg till bokm�rken|L�gg till aktuell fj�rrkatalog som bokm�rke
ImageIndex6ShortCutB@  TActionConsoleActionTagCategoryCommandCaption�ppna &terminalf�nsterHelpKeyword
ui_consoleHint��ppna terminalf�nster|�ppnar terminalf�nster som till�ter k�rande av godtyckligt extrakommando (med undantag av de som kr�ver anv�ndarinput)
ImageIndex7ShortCutT@  TActionPuttyActionTagCategoryCommandCaption�ppna session i &PuTTYHelpKeyword0integration_app#opening_current_session_in_puttyHintX�ppna session i PuTTY|Starta PuTTY SSH-terminalprogram och �ppna aktuell session med den
ImageIndex@ShortCutP@  TActionLocalExploreDirectoryActionTagCategoryLocal DirectoryCaption&Utforska katalogHint*�ppnar utforskaren i aktuell lokal katalog
ImageIndex8ShortCutE�    TActionCurrentOpenActionTagCategoryFocused OperationCaption&�ppnaHelpKeyword	task_editHintN�ppna dokument|�ppnar valt dokument med program som filtypen �r associerad med
ImageIndex:  TActionSynchronizeBrowsingActionTagCategoryCommand	AutoCheck	CaptionSynkronisera &bl�ddringHelpKeyword"task_navigate#synchronize_browsingHintGSynkronisera bl�ddring|Synkronisera lokal och fj�rrkatalogens bl�ddring
ImageIndex;ShortCutB�    TActionAddEditLinkActionTagCategoryCommandCaptionL�gg till/redigera &l�nk...HelpKeyword	task_linkHintSL�gg till/redigera l�nk|L�gger till ny l�nk/genv�g eller redigerar vald l�nk/genv�g
ImageIndex<  TActionAddEditLinkContextActionTagCategoryCommandCaptionRedigera &l�nk...HelpKeyword	task_linkHint'Redigera l�nk|Redigera vald l�nk/genv�g
ImageIndex<  TActionCloseApplicationActionTagCategory5Toolbar Operation (selected + rename + mkdir + close)Caption&AvslutaHintEAvsluta applikation|Avsluta �ppnade sessioner och st�ng applikationen
ImageIndex=  TActionOpenedSessionsActionTagCategorySessionCaption&�ppna sessionerHelpKeyword&task_connections#switching_connectionsHint-V�lj session|V�lj �ppnad session att aktivera
ImageIndex>  TActionDuplicateSessionActionTagCategorySessionCaption&Dubblera sessionHelpKeywordtask_connectionsHintaDubblera session|�ppnar samma session igen (h�ll nere SHIFT f�r att �ppna den i ett nytt f�nster)
ImageIndex[  TActionNewLinkActionTagCategoryCommandCaption&L�nk...HelpKeyword	task_linkHintSkapa l�nl|Skapa ny l�nk/genv�g
ImageIndex<  TActionCustomCommandsActionTagCategoryCommandCaptionEgna &kommandonHelpKeywordremote_command#custom_commandsHint+K�r egna kommandon med de markerade filerna  TActionCustomCommandsCustomizeActionTagCategoryCommandCaption&Anpassa...HelpKeywordui_pref_commandsHintAnpassa egna kommandon
ImageIndex  TActionCustomCommandsEnterActionTagCategoryCommandCaptionL�&gg in...HelpKeyword8remote_command#executing_and_configuring_custom_commandsHint!L�gg in egna kommandon f�r ad hoc
ImageIndexZ  TAction CustomCommandsEnterFocusedActionTagCategoryCommandCaptionL�&gg in...HelpKeyword8remote_command#executing_and_configuring_custom_commandsHint!L�gg in egna kommandon f�r ad hoc
ImageIndexZ  TActionCheckForUpdatesActionTagCategoryHelpCaptionS�k efter &uppdateringarHelpKeywordupdatesHint/Fr�gar applikationens webbsida om uppdateringar
ImageIndex?  TActionDonatePageActionTagCategoryHelpCaption&DoneraHintC�ppnar webbl�saren och g�r till programmets webbsida f�r donationer  TActionCustomCommandsLastActionTagCategoryCommandCaptionCustomCommandsLastActionHelpKeyword8remote_command#executing_and_configuring_custom_commands  TActionCustomCommandsLastFocusedActionTagCategoryCommandCaptionCustomCommandsLastFocusedActionHelpKeyword8remote_command#executing_and_configuring_custom_commands  TActionFileSystemInfoActionTagCategoryCommandCaption&Server/protokollinformationHelpKeyword	ui_fsinfoHint Visa server/protokollinformation
ImageIndex  TActionClearCachesActionTagCategoryCommandCaption&Rensa cacheHelpKeyworddirectory_cacheHint0Rensa cache f�r kataloglistning och katalogbyten  TActionFullSynchronizeActionTagCategoryCommandCaption&Synkronisera...HelpKeywordtask_synchronize_fullHint+Synkronisera lokal katalog med fj�rrkatalog
ImageIndexBShortCutS@  TActionRemoteMoveToFocusedActionTagCategoryFocused OperationCaption&Flytta till...HelpKeyword'task_move_duplicate#moving_remote_filesHint/Flytta|Flytta markerade filer till fj�rrkatalog  TActionShowHiddenFilesActionTagCategoryViewCaptionVisa/&d�lj d&olda filerHelpKeywordui_file_panel#special_filesHint(V�xla visning av dolda filer i panel(er)ShortCutH�    TActionLocalPathToClipboardActionTagCategoryLocal DirectoryCaptionKopiera s&�kv�g till urklippHelpKeyword#filenames#current_working_directoryHint)Kopiera aktuell lokal s�kv�g till urklipp  TActionRemotePathToClipboardActionTagCategoryRemote DirectoryCaptionKopiera s&�kv�g till urklippHelpKeyword#filenames#current_working_directoryHint(Kopiera aktuell fj�rrs�kv�g till urklipp  TActionFileListToCommandLineActionTagCategorySelected OperationCaptionIn&foga till kommandoradHelpKeywordfilenames#command_lineHint/Infoga markerade filers namn till kommandoradenShortCut@  TActionFileListToClipboardActionTagCategorySelected OperationCaption&Kopiera till urklippHelpKeywordfilenames#file_nameHint*Kopiera markerade filers namn till urklippShortCutC`  TActionFullFileListToClipboardActionTagCategorySelected OperationCaption*Kopiera till urklipp (inklusive s&�kv�gar)HelpKeywordfilenames#file_nameHint;Kopiera markerade filers namn inklusive s�kv�g till urklippShortCutC�    TActionQueueGoToActionTagCategoryQueueCaption&G� tillHelpKeywordui_queue#managing_the_queueHintG� till �verf�ringsk�listan
ImageIndexJShortCutQ@  TActionQueueItemUpActionTagCategoryQueueCaptionFlytta &uppHelpKeywordui_queue#managing_the_queueHint/Flytta upp vald k�post f�r att utf�ras tidigare
ImageIndexH  TActionQueueItemDownActionTagCategoryQueueCaptionFlytta &nerHelpKeywordui_queue#managing_the_queueHint-Flytta ner vald k�post f�r att utf�ras senare
ImageIndexI  TActionQueueToggleShowActionTagCategoryQueueCaption&K�HintVisa/d�lj k�lista
ImageIndexJ  TActionQueueShowActionTagCategoryQueueCaptionVi&saHelpKeywordui_queueHintVisa k�lista  TActionQueueHideWhenEmptyActionTagCategoryQueueCaptionD�lj ifall &tomHelpKeywordui_queueHintD�lj k�listan n�r den �r tom  TActionQueueHideActionTagCategoryQueueCaption&D�ljHelpKeywordui_queueHintD�lj k�lista  TActionQueueToolbarActionTagCategoryQueueCaption&Verktygsf�ltHint:D�lj/visa verktygsf�ltet f�r k�listan (p� k�listans panel)  TActionQueuePreferencesActionTagCategoryQueueCaptionA&npassa...HelpKeywordui_pref_backgroundHintAnpassa k�lista
ImageIndex  TActionPasteActionTagCategoryCommandCaptionK&listra inHelpKeyword task_upload#using_copy_amp:pasteHint@Klistra in filer fr�n urklipp till aktuell katalog i aktiv panel
ImageIndexKShortCutV@  TActionNewFileActionTagCategoryCommandCaption&Fil...HelpKeyword	task_editHint0Skapa fil|Skapar ny fil och �ppnas den i editorn
ImageIndexM  TActionEditorListCustomizeActionTagCategoryCommandCaption&Konfigurera...HelpKeywordui_pref_editorHintSkr�ddarsy editorer
ImageIndex  TActionRemoteCopyToFocusedActionTagCategoryFocused OperationCaption&Dubblera...HelpKeyword,task_move_duplicate#duplicating_remote_filesHint2Dubblera|Dubbleras valda filer till fj�rrkatalogen
ImageIndexN  TActionRemoteCopyToActionTagCategorySelected OperationCaption&Dubblera...HelpKeyword,task_move_duplicate#duplicating_remote_filesHint1Dubblera|Dubblera valda filer till fj�rrkatalogen
ImageIndexN  TActionUrlToClipboardActionTagCategorySelected OperationCaptionKopiera &URL till urklippHelpKeywordfilenames#file_urlHint*Kopiera URL'er av valda filer till urklipp  TActionTableOfContentsActionTagCategoryHelpCaption	I&nneh�llHintD�ppnar webbl�sare och g�r till dokumentationens inneh�llsf�rteckning
ImageIndexOShortCutp  TActionFileListFromClipboardActionTagCategorySelected OperationCaption&Transfer Files in ClipboardHint+Transfer files whose names are in clipboard  TActionRemoteCopyActionTagCategorySelected OperationCaptionLadda &ner...HelpKeywordtask_downloadHint Ladda ner|Ladda ner vald fil(er)
ImageIndexY  TActionLocalCopyActionTagCategorySelected OperationCaptionLadda &upp...HelpKeywordtask_uploadHint Ladda upp|Ladda upp vald fil(er)
ImageIndexX  TActionCurrentDeleteAlternativeActionTagCategorySelected OperationCaption&Ta bortHelpKeywordtask_deleteHintTa bort|Ta bort vald fil(er)
ImageIndex  TActionCurrentEditAlternativeActionTagCategorySelected OperationCaption&Redigera (alternativ)HelpKeyword	task_editHint=Redigera (alternativ)|Redigera vald fil med alternativ editor  TActionCurrentEditWithActionTagCategorySelected OperationCaptionRedigera &med...HelpKeyword	task_editHint:Redigera med|Redigera vald fil(er) med editorn som ni valt  TActionDownloadPageActionTagCategoryHelpCaption
Ladda &nerHint>�ppnar webbl�sare och g�r till applikationens nerladdningssida  TActionUpdatesPreferencesActionTagCategoryHelpCaptionKonfi&gurera...HelpKeywordui_pref_updatesHintBKonfigurera automatisk kontroll av uppdateringar f�r applikationen
ImageIndex  TActionShowUpdatesActionTagCategoryHelpCaption&Visa uppdateringarHelpKeywordupdatesHint�Visa information om applikationens uppdateringar|Visa information om applikationens uppdateringar (f�rfr�gar applikationens hemsida om informationen inte �r tillg�nglig vid tidpunkten)
ImageIndexQ  TActionPresetsPreferencesActionTagCategoryViewCaption&Konfigurera...HelpKeywordui_pref_presetsHint-Konfigurera f�rinst�llningar f�r �verf�ringar
ImageIndex  TActionLockToolbarsActionTagCategoryViewCaption&L�s verktygsf�ltHelpKeywordui_toolbarsHint2Hindra flyttning och dockning av alla verktygsf�lt  TActionCustomCommandsBandActionTagCategoryViewCaptionEgna ko&mmandoknapparHelpKeywordui_toolbarsHint)D�lj/visa verktygsf�lt f�r egna kommandon  TActionColorMenuActionTagCategoryViewCaptionF&�rgHelpKeywordtask_connections#session_colorHint�ndra f�rg p� aktuell session  TActionColorDefaultActionTagCategoryViewCaption	&StandardHelpKeywordtask_connections#session_colorHint2�terst�ll session (panel) f�rg till systemstandard  TActionColorPickActionTagCategoryViewCaptionFl%er f�rger...HelpKeywordtask_connections#session_colorHintV�lj f�rg p� session (panel)  TActionAutoReadDirectoryAfterOpActionTagCategoryViewCaptionLadda auto&matisk om katalogHint;�ndra automatisk omladdning av fj�rrkatalog efter operationShortCutR�    TActionQueueItemPauseActionTagCategoryQueueCaption&PausaHelpKeywordui_queue#managing_the_queueHintPausa vald k�post
ImageIndexS  TActionQueueItemResumeActionTagCategoryQueueCaption
&�terupptaHelpKeywordui_queue#managing_the_queueHint�teruppta vald pausad k�post
ImageIndexF  TActionQueuePauseAllActionTagCategoryQueueCaption&Pausa allaHelpKeywordui_queue#managing_the_queueHintPausa alla k�poster som k�rs
ImageIndexT  TActionQueueResumeAllActionTagCategoryQueueCaption&�teruppta allaHelpKeywordui_queue#managing_the_queueHint�teruppta alla pausade k�poster
ImageIndexU  TActionQueueDisconnectOnceEmptyActionTagCategoryQueueCaptionKo&ppla ifr�n ifall tomHelpKeywordui_queueHint#Koppla ifr�n session n�r k�n �r tom
ImageIndexW  TActionRestoreSelectionActionTagCategory	SelectionCaption&�terst�ll markeringHelpKeywordui_file_panel#selecting_filesHint�terst�ll f�reg�ende markering
ImageIndexV  TActionCurrentEditFocusedActionTagCategoryFocused OperationCaption	&RedigeraHelpKeyword	task_editHintRedigera|Redigera vald fil(er)
ImageIndex9  TActionNewDirActionTagCategoryCommandCaptionKatalo&g...HelpKeywordtask_create_directoryHintSkapa katalog|Skapa ny katalog
ImageIndex  TActionQueueShutDownOnceEmptyActionTagCategoryQueueCaption&Str�ng av datornHelpKeywordui_queueHintStr�ng av datorn n�r k�n �r tom
ImageIndex]  TActionQueueIdleOnceEmptyActionTagCategoryQueueCaption&F�rbli idleChecked	HelpKeywordui_queueHintF�rbli idle n�r k�n �r tom
ImageIndex^  TActionQueueCycleOnceEmptyActionTagCategoryQueueCaption&Tom k�HelpKeywordui_queueHint*�ndra �tg�rd som ska utf�ras d� k�n �r tom
ImageIndex^  TTBEditActionQueueItemSpeedActionTagCategoryQueueHelpKeywordui_queue#managing_the_queueHint%�ndra hastighetsgr�ns f�r vald k�postEditCaption
&Hastighet  TActionLocalFilterActionTag	CategoryLocal DirectoryCaption&Filtrera...HelpKeywordui_file_panel#filterHintFiltrera|Filtrera visade filer
ImageIndex\  TActionRemoteFilterActionTagCategoryRemote DirectoryCaption
&Filter...HelpKeywordui_file_panel#filterHintFilter|Filtrera visade filer
ImageIndex\  TActionFindFilesActionTagCategoryCommandCaptionS�&k filer..HelpKeyword	task_findHint!S�k filer|S�k filer och kataloger
ImageIndex_   TTBXPopupMenuExplorerBarPopupImagesGlyphsModule.ExplorerImagesLeft� TopP TTBXItemAddress2ActionExplorerAddressBandAction  TTBXItemStandardButtons1ActionExplorerToolbarBandAction  TTBXItemSelectionButtons1ActionExplorerSelectionBandAction  TTBXItemSessionButtons2ActionExplorerSessionBandAction  TTBXItemPreferencesButtons1ActionExplorerPreferencesBandAction  TTBXItemSortButtons3ActionExplorerSortBandAction  TTBXItemTBXItem3ActionExplorerUpdatesBandAction  TTBXItemTBXItem4ActionExplorerTransferBandAction  TTBXItem	TBXItem16Action ExplorerCustomCommandsBandAction  TTBXItemTBXItem7ActionLockToolbarsAction  TTBXSeparatorItemN5  TTBXItem
StatusBar2ActionStatusBarAction  TTBXSeparatorItemN72  TTBXSubmenuItemQueue7Caption&K�HelpKeywordui_queueHintKonfigurera k�lista TTBXItemShow6ActionQueueShowAction	RadioItem	  TTBXItemHidewhenEmpty6ActionQueueHideWhenEmptyAction	RadioItem	  TTBXItemHide5ActionQueueHideAction	RadioItem	  TTBXSeparatorItemN71  TTBXItemToolbar5ActionQueueToolbarAction  TTBXSeparatorItemN70  TTBXItem
Customize5ActionQueuePreferencesAction   TTBXItemTree4ActionRemoteTreeAction   TTimerSessionIdleTimerEnabledInterval�OnTimerSessionIdleTimerTimerLeft TopP  TTBXPopupMenuCommanderBarPopupImagesGlyphsModule.ExplorerImagesLeft�Top TTBXItemStandardButtons3ActionCommanderToolbarBandAction  TTBXItemSessionButtons5ActionCommanderSessionBandAction  TTBXItemSelectionButtons3ActionCommanderSelectionBandAction  TTBXItemPreferencesButtons4ActionCommanderPreferencesBandAction  TTBXItemSortButtons2ActionCommanderSortBandAction  TTBXItemCommandsButtons2ActionCommanderCommandsBandAction  TTBXItemTBXItem2ActionCommanderUpdatesBandAction  TTBXItemTBXItem5ActionCommanderTransferBandAction  TTBXItem	TBXItem14Action!CommanderUploadDownloadBandAction  TTBXItem	TBXItem15Action!CommanderCustomCommandsBandAction  TTBXItemTBXItem6ActionLockToolbarsAction  TTBXSeparatorItemN26  TTBXItemCommandLine2ActionCommandLinePanelAction  TTBXItemCommandsToolbar1ActionToolBarAction  TTBXItem
StatusBar8ActionStatusBarAction  TTBXSeparatorItemN27  TTBXSubmenuItemLocalPanel1Caption&Lokal panelHelpKeywordui_file_panelHint"�ndra den lokala panelens utseende TTBXItemHistoryButtons3ActionCommanderLocalHistoryBandAction  TTBXItemNavigationButtons3Action"CommanderLocalNavigationBandAction  TTBXSeparatorItemN23  TTBXItemTree7ActionLocalTreeAction  TTBXSeparatorItemN77  TTBXItem
StatusBar6ActionLocalStatusBarAction   TTBXSubmenuItemRemotePanel2Caption&Fj�rrpanelHelpKeywordui_file_panelHint�ndra fj�rrpanelens utseende TTBXItemHistoryButtons4Action CommanderRemoteHistoryBandAction  TTBXItemNavigationButtons4Action#CommanderRemoteNavigationBandAction  TTBXSeparatorItemN25  TTBXItemTree8ActionRemoteTreeAction  TTBXSeparatorItemN78  TTBXItem
StatusBar7ActionRemoteStatusBarAction   TTBXSubmenuItemOptions1Caption&K�HelpKeywordui_queueHintKonfigurera k�lista TTBXItemShow5ActionQueueShowAction	RadioItem	  TTBXItemHidewhenEmpty5ActionQueueHideWhenEmptyAction	RadioItem	  TTBXItemHide4ActionQueueHideAction	RadioItem	  TTBXSeparatorItemN69  TTBXItemToolbar4ActionQueueToolbarAction  TTBXSeparatorItemN68  TTBXItem
Customize4ActionQueuePreferencesAction    TTBXPopupMenuRemotePanelPopupImagesGlyphsModule.ExplorerImagesLeft8Top TTBXItem	TBXItem32ActionRemoteRefreshAction  TTBXItem	TBXItem30ActionRemoteAddBookmarkAction  TTBXItemCopyPathtoClipboard1ActionRemotePathToClipboardAction  TTBXItemOpenDirectoryBookmark1ActionRemoteOpenDirAction  TTBXItem	TBXItem26ActionRemoteFilterAction  TTBXSeparatorItemN51  TTBXItemHistoryButtons5Action CommanderRemoteHistoryBandAction  TTBXItemNavigationButtons5Action#CommanderRemoteNavigationBandAction  TTBXSeparatorItemN28  TTBXItemTree5ActionRemoteTreeAction  TTBXSeparatorItemN75  TTBXItem
StatusBar9ActionRemoteStatusBarAction   TTBXPopupMenuLocalPanelPopupImagesGlyphsModule.ExplorerImagesLeft8TopP TTBXItem	TBXItem34ActionLocalRefreshAction  TTBXItem	TBXItem31ActionLocalAddBookmarkAction  TTBXItemCopyPathtoClipboard2ActionLocalPathToClipboardAction  TTBXItemOpenDirectoryBookmark2ActionLocalOpenDirAction  TTBXItem	TBXItem27ActionLocalFilterAction  TTBXSeparatorItemN52  TTBXItemHistoryButtons6ActionCommanderLocalHistoryBandAction  TTBXItemNavigationButtons6Action"CommanderLocalNavigationBandAction  TTBXSeparatorItemN29  TTBXItemTree6ActionLocalTreeAction  TTBXSeparatorItemN76  TTBXItemStatusBar10ActionLocalStatusBarAction   TTBXPopupMenuLocalDirViewColumnPopupImagesGlyphsModule.ExplorerImagesLeft� TopX TTBXItemSortAscending1ActionSortColumnAscendingAction  TTBXItemSortDescending1ActionSortColumnDescendingAction  TTBXItemLocalSortByExtColumnPopupItemActionLocalSortByExtAction  TTBXItemHidecolumn1ActionHideColumnAction  TTBXSeparatorItemN37  TTBXSubmenuItemShowcolumns3CaptionVisa &kolumnerHelpKeywordui_file_panel#selecting_columnsHint%V�lj kolumner som ska visas i panelen TTBXItemName3ActionShowHideLocalNameColumnAction  TTBXItemSize3ActionShowHideLocalSizeColumnAction  TTBXItemType2ActionShowHideLocalTypeColumnAction  TTBXItemModification3Action ShowHideLocalChangedColumnAction  TTBXItemAttributes3ActionShowHideLocalAttrColumnAction    TTBXPopupMenuRemoteDirViewColumnPopupImagesGlyphsModule.ExplorerImagesLeft�TopX TTBXItem	MenuItem1ActionSortColumnAscendingAction	RadioItem	  TTBXItem	MenuItem2ActionSortColumnDescendingAction	RadioItem	  TTBXItemRemoteSortByExtColumnPopupItemActionRemoteSortByExtAction  TTBXItemHidecolumn2ActionHideColumnAction  TTBXSeparatorItemN38  TTBXSubmenuItemShowcolumns4CaptionVisa &kolumnerHelpKeywordui_file_panel#selecting_columnsHint%V�lj kolumner som ska visas i panelen TTBXItemName4ActionShowHideRemoteNameColumnAction  TTBXItemSize4ActionShowHideRemoteSizeColumnAction  TTBXItemTBXItem8ActionShowHideRemoteTypeColumnAction  TTBXItemModification4Action!ShowHideRemoteChangedColumnAction  TTBXItemPermissions1Action ShowHideRemoteRightsColumnAction  TTBXItemOwner2ActionShowHideRemoteOwnerColumnAction  TTBXItemGroup2ActionShowHideRemoteGroupColumnAction  TTBXItemTBXItem1Action$ShowHideRemoteLinkTargetColumnAction    TTBXPopupMenu
QueuePopupImagesGlyphsModule.ExplorerImagesOnPopupQueuePopupPopupLeft�Top�  TTBXItem
ShowQuery1ActionQueueItemQueryAction  TTBXItem
ShowError1ActionQueueItemErrorAction  TTBXItemShowPrompt1ActionQueueItemPromptAction  TTBXSeparatorItemN53  TTBXItemExecuteNow1ActionQueueItemExecuteAction  TTBXItemTBXItem9ActionQueueItemPauseAction  TTBXItem	TBXItem10ActionQueueItemResumeAction  TTBXItemDelete4ActionQueueItemDeleteAction  TTBXComboBoxItemQueuePopupSpeedComboBoxItemActionQueueItemSpeedAction  TTBXSeparatorItemN54  TTBXItemMoveUp1ActionQueueItemUpAction  TTBXItem	MoveDown1ActionQueueItemDownAction  TTBXSeparatorItemN67  TTBXSubmenuItemTBXSubmenuItem1Caption&AllaHelpKeywordui_queue#managing_the_queueHint$Administrationskommandon f�r k�massa TTBXItem	TBXItem11ActionQueuePauseAllAction  TTBXItem	TBXItem12ActionQueueResumeAllAction   TTBXSubmenuItemTBXSubmenuItem3ActionQueueCycleOnceEmptyActionDropdownCombo	 TTBXItem	TBXItem28ActionQueueIdleOnceEmptyAction	RadioItem	  TTBXItem	TBXItem13ActionQueueDisconnectOnceEmptyAction	RadioItem	  TTBXItem	TBXItem29ActionQueueShutDownOnceEmptyAction	RadioItem	   TTBXSubmenuItemQueue2Caption&AlternativHelpKeywordui_queueHintKonfigurera k�lista TTBXItemShow4ActionQueueShowAction	RadioItem	  TTBXItemHidewhenEmpty4ActionQueueHideWhenEmptyAction	RadioItem	  TTBXItemHide3ActionQueueHideAction	RadioItem	  TTBXSeparatorItemN66  TTBXItemToolbar3ActionQueueToolbarAction  TTBXSeparatorItemN65  TTBXItem
Customize3ActionQueuePreferencesAction    TTBXPopupMenuRemoteDirViewPopupImagesGlyphsModule.ExplorerImagesLefthTop� TTBXSubmenuItemGoTo4Caption&G� tillHelpKeywordtask_navigateHintG� till katalog TTBXItemOpenDirectoryBookmark3ActionRemoteOpenDirAction  TTBXSeparatorItemN81  TTBXItemParentDirectory4ActionRemoteParentDirAction  TTBXItemRootDirectory4ActionRemoteRootDirAction  TTBXItemHomeDirectory4ActionRemoteHomeDirAction  TTBXSeparatorItemN80  TTBXItemBack4ActionRemoteBackAction  TTBXItemForward4ActionRemoteForwardAction   TTBXItemRefresh4ActionRemoteRefreshAction  TTBXItemAddToBookmarks4ActionRemoteAddBookmarkAction  TTBXItemCopyPathtoClipboard6ActionRemotePathToClipboardAction  TTBXSeparatorItemN79  TTBXSubmenuItemTBXSubmenuItem26Caption&NyHelpKeyword
task_indexHintSkapa objekt|Skapa nytt objekt TTBXItem
TBXItem135ActionNewFileAction  TTBXItem
TBXItem136ActionNewDirAction  TTBXItem
TBXItem209ActionNewLinkAction    TTBXPopupMenuLocalDirViewPopupImagesGlyphsModule.ExplorerImagesLeft�Top� TTBXSubmenuItemGoTo5Caption&G� tillHelpKeywordtask_navigateHintG� till katalog TTBXItemOpenDirectoryBookmark4ActionLocalOpenDirAction  TTBXItemExploreDirectory2ActionLocalExploreDirectoryAction  TTBXSeparatorItemN84  TTBXItemParentDirectory5ActionLocalParentDirAction  TTBXItemRootDirectory5ActionLocalRootDirAction  TTBXItemHomeDirectory5ActionLocalHomeDirAction  TTBXSeparatorItemN83  TTBXItemBack5ActionLocalBackAction  TTBXItemForward5ActionLocalForwardAction   TTBXItemRefresh5ActionLocalRefreshAction  TTBXItemAddToBookmarks5ActionLocalAddBookmarkAction  TTBXItemCopyPathtoClipboard7ActionLocalPathToClipboardAction  TTBXSeparatorItemN82  TTBXItemCreateDirectory4ActionCurrentCreateDirAction   TTBXPopupMenuRemoteAddressPopupImagesGlyphsModule.ExplorerImagesLeft� Top� TTBXItem	TBXItem33ActionRemoteRefreshAction  TTBXItem	TBXItem24ActionRemoteAddBookmarkAction  TTBXItem	TBXItem25ActionRemotePathToClipboardAction  TTBXSeparatorItemTBXSeparatorItem1  TTBXItem	TBXItem17ActionRemoteOpenDirAction  TTBXSubmenuItemTBXSubmenuItem2Caption&G� tillHelpKeywordtask_navigateHintG� till katalog TTBXItem	TBXItem18ActionRemoteParentDirAction  TTBXItem	TBXItem19ActionRemoteRootDirAction  TTBXItem	TBXItem20ActionRemoteHomeDirAction  TTBXSeparatorItemTBXSeparatorItem2  TTBXItem	TBXItem21ActionRemoteBackAction  TTBXItem	TBXItem22ActionRemoteForwardAction        TPF0TOpenDirectoryDialogOpenDirectoryDialogLeft�Top� HelpType	htKeywordHelpKeyword
ui_opendirBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionOpen directoryClientHeightNClientWidth�Color	clBtnFace
ParentFont	OldCreateOrder	PositionpoMainFormCenterOnShowFormShow
DesignSize�N PixelsPerInch`
TextHeight TLabel	EditLabelLeftTopWidthHHeightCaption&�ppna katalog:  TIEComboBoxLocalDirectoryEditLeftTopWidth4HeightAnchorsakLeftakTopakRight 
ItemHeightTabOrderTextLocalDirectoryEditOnChangeDirectoryEditChange  TIEComboBoxRemoteDirectoryEditLeftTopWidth�HeightAnchorsakLeftakTopakRight 
ItemHeight	MaxLength�TabOrder TextRemoteDirectoryEditOnChangeDirectoryEditChange  TButtonOKBtnLeft� Top,WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeft� Top,WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TPageControlPageControlLeftTop8Width�Height� 
ActivePageSessionBookmarksSheetAnchorsakLeftakTopakRightakBottom TabIndex TabOrder 	TTabSheetSessionBookmarksSheetTagCaptionSessionsbokm�rken
DesignSizez�   TListBoxSessionBookmarksListTagLeft
Top	WidthHeight� AnchorsakLeftakTopakRightakBottom DragModedmAutomatic
ItemHeightTabOrder OnClickBookmarksListClick
OnDblClickBookmarksListDblClick
OnDragDropBookmarksListDragDrop
OnDragOverBookmarksListDragOver	OnEndDragBookmarksListEndDrag	OnKeyDownBookmarksListKeyDownOnStartDragBookmarksListStartDrag  TButtonAddSessionBookmarkButtonTagLeftTop	WidthSHeightAnchorsakTopakRight Caption
&L�gg tillTabOrderOnClickAddBookmarkButtonClick  TButtonRemoveSessionBookmarkButtonTagLeftTop)WidthSHeightAnchorsakTopakRight Caption&Ta bortTabOrderOnClickRemoveBookmarkButtonClick  TButtonUpSessionBookmarkButtonTag�LeftTop� WidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickBookmarkButtonClick  TButtonDownSessionBookmarkButtonTagLeftTop� WidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickBookmarkButtonClick   	TTabSheetSharedBookmarksSheetTagCaptionDelade bokm�rken
ImageIndex
DesignSizez�   TListBoxSharedBookmarksListTagLeft
Top	WidthHeight� AnchorsakLeftakTopakRightakBottom DragModedmAutomatic
ItemHeightTabOrder OnClickBookmarksListClick
OnDblClickBookmarksListDblClick
OnDragDropBookmarksListDragDrop
OnDragOverBookmarksListDragOver	OnEndDragBookmarksListEndDrag	OnKeyDownBookmarksListKeyDownOnStartDragBookmarksListStartDrag  TButtonAddSharedBookmarkButtonTagLeftTop	WidthSHeightAnchorsakTopakRight Caption
&L�gg tillTabOrderOnClickAddBookmarkButtonClick  TButtonRemoveSharedBookmarkButtonTagLeftTop)WidthSHeightAnchorsakTopakRight Caption&Ta bortTabOrderOnClickRemoveBookmarkButtonClick  TButtonUpSharedBookmarkButtonTag�LeftTop� WidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickBookmarkButtonClick  TButtonDownSharedBookmarkButtonTagLeftTop� WidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickBookmarkButtonClick  TButtonShortCutSharedBookmarkButtonTagLeftTopIWidthSHeightAnchorsakTopakRight Caption
&Genv�g...TabOrderOnClickShortCutBookmarkButtonClick    TButtonLocalDirectoryBrowseButtonLeft@TopWidthKHeightAnchorsakTopakRight CaptionBl�dd&ra...TabOrderOnClickLocalDirectoryBrowseButtonClick  TButtonSwitchButtonLeftTop,WidthyHeightAnchorsakLeftakBottom CaptionP&latsprofiler...ModalResultTabOrderOnClickSwitchButtonClick  TButton
HelpButtonLeft@Top,WidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrderOnClickHelpButtonClick    TPF0TPreferencesDialogPreferencesDialogLeft�Top� HelpType	htKeywordHelpKeywordui_preferencesBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionInst�llningarClientHeight�ClientWidthColor	clBtnFace
ParentFont	OldCreateOrder	PositionpoMainFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize� PixelsPerInch`
TextHeight TButtonOKButtonLeft� TopqWidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCloseButtonLeftRTopqWidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TPanel	MainPanelLeft Top WidthHeightkAlignalTopAnchorsakLeftakTopakRightakBottom 
BevelOuterbvNoneTabOrder  TPageControlPageControlLeft� Top Width}Heightk
ActivePagePreferencesSheetAlignalClient	MultiLine	Style	tsButtonsTabOrderTabStopOnChangePageControlChange 	TTabSheetPreferencesSheetTagHintMilj�HelpType	htKeywordHelpKeywordui_pref_environmentCaptionGen
ImageIndex
TabVisible
DesignSizeua  	TGroupBoxCommonPreferencesGroupLeftTopWidtheHeight AnchorsakLeftakTopakRight CaptionBekr�ftelserTabOrder 
DesignSizee   	TCheckBoxConfirmOverwritingCheckLeftTop,WidthEHeightAnchorsakLeftakTopakRight Caption&�verskrivning av filerTabOrderOnClickControlChange  	TCheckBoxConfirmDeletingCheckLeftTopCWidthEHeightAnchorsakLeftakTopakRight Caption%&Borttagning av filer (rekommenderad)TabOrderOnClickControlChange  	TCheckBoxConfirmClosingSessionCheckLeftTop� WidthEHeightAnchorsakLeftakTopakRight CaptionA&vsluta applikationenTabOrderOnClickControlChange  	TCheckBoxDDTransferConfirmationCheckLeftTop� WidthEHeightAnchorsakLeftakTopakRight CaptionD&ra && sl�pp-operationerTabOrderOnClickControlChange  	TCheckBoxContinueOnErrorCheckLeftTop� WidthEHeightAnchorsakLeftakTopakRight Caption(Forts�tt vid &fel (avancerade anv�ndare)TabOrder	OnClickControlChange  	TCheckBoxConfirmExitOnCompletionCheckLeftTop� WidthEHeightAnchorsakLeftakTopakRight Caption-Avsluta a&pplikationen vid slutf�rd operationTabOrderOnClickControlChange  	TCheckBoxConfirmResumeCheckLeftTopqWidthEHeightAnchorsakLeftakTopakRight Caption&�teruppta �verf�ringTabOrderOnClickControlChange  	TCheckBoxConfirmCommandSessionCheckLeftTop� WidthEHeightAnchorsakLeftakTopakRight Caption�ppna separat &skalsessionTabOrderOnClickControlChange  	TCheckBoxConfirmRecyclingCheckLeftTopZWidthEHeightAnchorsakLeftakTopakRight Caption &Flytta filer till papperskorgenTabOrderOnClickControlChange  	TCheckBoxConfirmTransferringCheckLeftTopWidthEHeightAnchorsakLeftakTopakRight Caption&�verf�ring av filerTabOrder OnClickControlChange   	TGroupBoxNotificationsGroupLeftTopWidtheHeightIAnchorsakLeftakTopakRight CaptionMeddelandenTabOrder
DesignSizeeI  TLabelBeepOnFinishAfterTextLeftXTopWidthHeightCaptions  	TCheckBoxBeepOnFinishCheckLeftTopWidthHeightAnchorsakLeftakTopakRight Caption8S&ystemljud n�r operationen �r klar, om den p�g�r mer �nTabOrder OnClickControlChange  TUpDownEditBeepOnFinishAfterEditLeftTopWidth9Height	AlignmenttaRightJustify	IncrementMaxValue�	MaxLengthTabOrderOnChangeControlChange  	TCheckBoxBalloonNotificationsCheckLeftTop.Width5HeightAnchorsakLeftakTopakRight CaptionHVisa ballong&meddelanden i aktivitetsf�ltets statusomr�de (systemf�ltet)TabOrderOnClickControlChange    	TTabSheetLogSheetTagHintLoggningHelpType	htKeywordHelpKeywordui_pref_loggingCaptionLog
ImageIndex
TabVisible
DesignSizeua  �TLoggingFrameLoggingFrameLeftTopWidthtHeightAnchorsakLeftakTopakRight TabOrder 
DesignSizet  �	TGroupBoxLoggingGroupWidthe
DesignSizee�   �TFilenameEditLogFileNameEdit2Width/  �TPanelLogFilePanelWidth1   �	TGroupBoxLogGroupWidthe    	TTabSheetGeneralSheetTagHint
Gr�nssnittHelpType	htKeywordHelpKeywordui_pref_interfaceCaptionInt
ImageIndex
TabVisible
DesignSizeua  TLabelLabel1LeftTop� WidthiHeight!AutoSizeCaptionWNotera: en �ndring i inst�llningen ger resultat f�rst vid n�sta uppstart av programmet.WordWrap	  �TGeneralSettingsFrameGeneralSettingsFrameLeftTopWidtheHeight� AnchorsakLeftakTopakRight TabOrder  �	TGroupBoxInterfaceGroupWidthj �TLabelCommanderDescriptionLabel2Width�   �TLabelExplorerDescriptionLabelWidth�     	TGroupBox
ThemeGroupLeftTop WidthiHeight4CaptionTemaTabOrder
DesignSizei4  TLabelLabel7LeftTopWidthMHeightCaptionGr�nssnitts&tema:FocusControl
ThemeCombo  	TComboBox
ThemeComboLeftxTopWidthqHeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrder Items.StringsSystem	Office XPOffice 2003     	TTabSheetPanelsSheetTagHintPanelerHelpType	htKeywordHelpKeywordui_pref_panelsCaptionPan
ImageIndex
TabVisible
DesignSizeua  	TGroupBoxPanelsRemoteDirectoryGroupLeftTop� WidtheHeightIAnchorsakLeftakTopakRight CaptionFj�rrkatalogTabOrder
DesignSizeeI  	TCheckBoxShowInaccesibleDirectoriesCheckLeftTopWidthEHeightAnchorsakLeftakTopakRight CaptionVis&a o�tkomliga katalogerTabOrder OnClickControlChange  	TCheckBoxAutoReadDirectoryAfterOpCheckLeftTop,WidthEHeightAnchorsakLeftakTopakRight Caption:Uppdatera auto&matisk katalog efter operation (CTRL+ALT+R)TabOrderOnClickControlChange   	TGroupBoxPanelsCommonGroupLeftTopWidtheHeight� AnchorsakLeftakTopakRight CaptionAllm�ntTabOrder 
DesignSizee�   	TCheckBoxShowHiddenFilesCheckLeftTopWidthEHeightAnchorsakLeftakTopakRight CaptionVi&sa dolda filer (CTRL+ALT+H)TabOrder OnClickControlChange  	TCheckBoxDefaultDirIsHomeCheckLeftTopCWidthEHeightAnchorsakLeftakTopakRight Caption Standardkatalog �r &hemkatalogenTabOrderOnClickControlChange  	TCheckBoxDeleteToRecycleBinCheckLeftTop,WidthEHeightAnchorsakLeftakTopakRight Caption'Ta bort lokala filer till papperskorgenTabOrderOnClickControlChange  	TCheckBoxPreservePanelStateCheckLeftTopZWidthEHeightAnchorsakLeftakTopakRight Caption0Kom i&h�g panelens' tillst�nd n�r session v�xlasTabOrderOnClickControlChange  	TCheckBoxRenameWholeNameCheckLeftTopqWidthEHeightAnchorsakLeftakTopakRight Caption#V�lj &hela namnet n�r filen d�ps omTabOrderOnClickControlChange   	TGroupBoxDoubleClickGroupLeftTop� WidtheHeightHAnchorsakLeftakTopakRight CaptionDubbelklickTabOrder
DesignSizeeH  TLabelDoubleClickActionLabelLeftTopWidth� HeightCaption&&Operation att utf�ra vid dubbelklick:FocusControlDoubleClickActionCombo  	TCheckBox"CopyOnDoubleClickConfirmationCheckLeft Top,Width4HeightAnchorsakLeftakTopakRight Caption*&Bekr�fta kopiera vid dubbelklickoperationTabOrderOnClickControlChange  	TComboBoxDoubleClickActionComboLeft� TopWidthlHeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrder OnChangeControlChangeItems.Strings�ppnaKopieraRedigera     	TTabSheetCommanderSheetTagHint	CommanderHelpType	htKeywordHelpKeywordui_pref_commanderCaptionCmd
ImageIndex
TabVisible
DesignSizeua  TLabelLabel3LeftTopWidthiHeightAnchorsakLeftakTopakRight AutoSizeCaptionPInst�llningar p� den h�r fliken g�ller endast f�r Norton Commander-gr�nssnittet.WordWrap	  	TGroupBoxPanelsGroupLeftTop&WidtheHeight� AnchorsakLeftakTopakRight CaptionPanelerTabOrder 
DesignSizee�   TLabelLabel8LeftTopWidthnHeightCaptionVal av &utforskarstil:FocusControlNortonLikeModeCombo  	TCheckBoxPreserveLocalDirectoryCheckLeftTop-WidthEHeightAnchorsakLeftakTopakRight Caption>&�ndra inte tillst�nd p� lokal paneler vid v�xlande av sessionTabOrderOnClickControlChange  	TCheckBoxSwappedPanelsCheckLeftTopEWidthEHeightAnchorsakLeftakTopakRight Caption3B&yt paneler (lokal till h�ger, fj�rr till v�nster)TabOrderOnClickControlChange  	TComboBoxNortonLikeModeComboLeft� TopWidth� HeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrder OnChangeControlChangeItems.StringsAldrigBara musMus och tangentbord   	TCheckBoxFullRowSelectCheckLeftTop]WidthEHeightAnchorsakLeftakTopakRight CaptionV�lja med h&ela radenTabOrderOnClickControlChange  	TCheckBoxTreeOnLeftCheckLeftTopuWidthEHeightAnchorsakLeftakTopakRight Caption&Visa &katalogtr�d v�nster om fillistanTabOrderOnClickControlChange   	TGroupBoxCommanderMiscGroupLeftTop� WidtheHeight5AnchorsakLeftakTopakRight Caption�vrigtTabOrder
DesignSizee5  	TCheckBoxUseLocationProfilesCheckLeftTopWidthEHeightAnchorsakLeftakTopakRight Caption3&Anv�nd platsprofiler ist�llet f�r katalogbokm�rkenTabOrder OnClickControlChange   	TGroupBoxCompareCriterionsGroupLeftTopWidtheHeightJAnchorsakLeftakTopakRight CaptionJ�mf�r katalogkriteriumTabOrder
DesignSizeeJ  	TCheckBoxCompareByTimeCheckLeftTopWidthEHeightAnchorsakLeftakTopakRight CaptionJ�mf�r efter &tidTabOrder OnClickControlChange  	TCheckBoxCompareBySizeCheckLeftTop-WidthEHeightAnchorsakLeftakTopakRight CaptionJ�mf�r efter &storlekTabOrderOnClickControlChange    	TTabSheetExplorerSheetTagHintUtforskarenHelpType	htKeywordHelpKeywordui_pref_explorerCaptionExp
ImageIndex
TabVisible
DesignSizeua  TLabelLabel4LeftTopWidthiHeightAnchorsakLeftakTopakRight AutoSizeCaptionGinst�llningar p� den h�r fliken g�ller endast f�r utforskargr�nssnittetWordWrap	  	TGroupBox	GroupBox2LeftTop&WidtheHeight6AnchorsakLeftakTopakRight CaptionVisaTabOrder 
DesignSizee6  	TCheckBoxShowFullAddressCheckLeftTopWidthEHeightAnchorsakLeftakTopakRight Caption.Vi&sa den fullst�ndiga s�kv�gen i adressf�ltetTabOrder OnClickControlChange    	TTabSheetTransferSheetTagHint
�verf�ringHelpType	htKeywordHelpKeywordui_pref_transferCaptionTran
ImageIndex
TabVisible �TCopyParamsFrameCopyParamsFrameLeft Top WidthHeightaHelpType	htKeyword
AutoScrollTabOrder    	TTabSheetEditorSheetTagHintEditorHelpType	htKeywordHelpKeywordui_pref_editorCaptionEdit
ImageIndex
TabVisible
DesignSizeua  	TGroupBoxInternalEditorGroupLeftTop� WidtheHeight� AnchorsakLeftakTopakRight CaptionAlternativ f�r intern editorTabOrder
DesignSizee�   TLabelEditorFontLabelLeft� TopWidth� HeightbAnchorsakLeftakTopakRight AutoSizeCaptionEditorFontLabelColor	clBtnFaceParentColor
OnDblClickEditorFontLabelDblClick  TLabelLabel9LeftTopOWidthEHeightCaption&Tabulatorstorlek:FocusControlEditorTabSizeEdit  TButtonEditorFontButtonLeftTopWidthiHeightAnchorsakTopakRight Caption&V�lj font...TabOrder OnClickEditorFontButtonClick  	TCheckBoxEditorWordWrapCheckLeftTop4Width~HeightAnchorsakLeftakTopakRight CaptionKo&rta av l�nga raderTabOrderOnClickControlChange  TUpDownEditEditorTabSizeEditLeftTop`WidthYHeight	AlignmenttaRightJustifyMaxValuecMinValueValue	MaxLengthTabOrderOnChangeControlChange   	TGroupBoxEditorPreferenceGroupLeftTopWidtheHeight� AnchorsakLeftakTopakRight CaptionEditorinst�llningarTabOrder 
DesignSizee�   	TListViewEditorListView2LeftTopWidthDHeight^AnchorsakLeftakTopakRightakBottom ColumnsCaptionMaskWidthF CaptionEditorWidth�  CaptionTextTagWidth-  ColumnClickDragModedmAutomaticHideSelection	OwnerData	ReadOnly		RowSelect	TabOrder 	ViewStylevsReportOnDataEditorListView2Data
OnDblClickEditorListView2DblClick	OnEndDragListViewEndDrag
OnDragDropEditorListView2DragDrop
OnDragOverListViewDragOver	OnKeyDownEditorListView2KeyDownOnSelectItemListViewSelectItemOnStartDragListViewStartDrag  TButtonAddEditorButtonLeftTop}WidthSHeightAnchorsakRightakBottom Caption&L�gg till...TabOrderOnClickAddEditEditorButtonClick  TButtonEditEditorButtonLeftpTop}WidthSHeightAnchorsakRightakBottom Caption&Redigera...TabOrderOnClickAddEditEditorButtonClick  TButtonUpEditorButtonLeftTop}WidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickUpDownEditorButtonClick  TButtonDownEditorButtonLeftTop� WidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickUpDownEditorButtonClick  TButtonRemoveEditorButtonLeftTop� WidthSHeightAnchorsakRightakBottom Caption&Ta bortTabOrderOnClickRemoveEditorButtonClick    	TTabSheetIntegrationSheetTag	HintIntegreringHelpType	htKeywordHelpKeywordui_pref_integrationCaptionInteg
ImageIndex
TabVisible
DesignSizeua  	TGroupBoxShellIconsGroupLeftTopWidtheHeight� AnchorsakLeftakTopakRight CaptionWindowsskalTabOrder 
DesignSizee�   TButtonDesktopIconButtonLeftTopWidthEHeightAnchorsakLeftakTopakRight CaptionSkapa en ikon p� skrivbor&detTabOrder OnClickIconButtonClick  TButtonQuickLaunchIconButtonLeftTop8WidthEHeightAnchorsakLeftakTopakRight CaptionSkapa en sna&bbstartsikonTabOrderOnClickIconButtonClick  TButtonSendToHookButtonLeftTopXWidthEHeightAnchorsakLeftakTopakRight Caption?Skapa genv�g f�r uppladdning i utforskarens '&Skicka till'-menyTabOrderOnClickIconButtonClick  TButtonRegisterAsUrlHandlerButtonLeftTop� WidthEHeightAnchorsakLeftakTopakRight Caption'Hantera adresser med scp:// och sftp://TabOrderOnClickRegisterAsUrlHandlerButtonClick  TButtonAddSearchPathButtonLeftTop� WidthEHeightAnchorsakLeftakTopakRight Caption0Addera s�kv�gen till WinSCP i milj�varibeln PATHTabOrderOnClickAddSearchPathButtonClick  TStaticTextShellIconsTextLeftToptWidthJHeightHint�F�r att l�gga till genv�gar, som �ppnar sparade sessioner direkt, anv�nd knappen 'Skalikon' p� ' sparade sessions' fliken i inloggningsdialogen	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption%Associera ikoner med sparde sessionerTabOrderTabStop	    	TTabSheetCustomCommandsSheetTag
Hint	KommandonHelpType	htKeywordHelpKeywordui_pref_commandsCaptionCmds
ImageIndex	
TabVisible
DesignSizeua  	TGroupBoxCustomCommandsGroupLeftTopWidtheHeightOAnchorsakLeftakTopakRightakBottom CaptionEgna kommandonTabOrder 
DesignSizeeO  	TListViewCustomCommandsViewLeftTopWidthDHeight� AnchorsakLeftakTopakRightakBottom ColumnsCaptionBeskrivningWidthU CaptionKommandoWidth�  CaptionL/FTagWidth# CaptionK/RTagWidth(  ColumnClickDragModedmAutomaticHideSelection	OwnerData	ReadOnly		RowSelect	TabOrder 	ViewStylevsReportOnDataCustomCommandsViewData
OnDblClickCustomCommandsViewDblClick	OnEndDragListViewEndDrag
OnDragDropCustomCommandsViewDragDrop
OnDragOverListViewDragOver	OnKeyDownCustomCommandsViewKeyDownOnSelectItemListViewSelectItemOnStartDragListViewStartDrag  TButtonAddCommandButtonLeftTopWidthSHeightAnchorsakRightakBottom Caption&L�gg till...TabOrderOnClickAddEditCommandButtonClick  TButtonRemoveCommandButtonLeftTop&WidthSHeightAnchorsakRightakBottom Caption&Ta bortTabOrderOnClickRemoveCommandButtonClick  TButtonUpCommandButtonLeftTopWidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickUpDownCommandButtonClick  TButtonDownCommandButtonLeftTop&WidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickUpDownCommandButtonClick  TButtonEditCommandButtonLeftpTopWidthSHeightAnchorsakRightakBottom Caption&Redigera...TabOrderOnClickAddEditCommandButtonClick    	TTabSheetDragDropSheetTagHintDra & sl�ppHelpType	htKeywordHelpKeywordui_pref_dragdropCaptionDragDrop
ImageIndex

TabVisible
DesignSizeua  	TGroupBoxDragDropDownloadsGroupLeftTopWidtheHeight� AnchorsakLeftakTopakRight CaptionDra && sl�pp nerladdningarTabOrder 
DesignSizee�   TLabelDDExtEnabledLabelLeft#TopDWidth9Height5AnchorsakLeftakTopakRight AutoSizeCaption�M�jligg�r direkt nerladdningar till vanliga lokala mappar (t. ex. utforskaren). Till�ter inte nerladdningar till andra destinationer (ZIP-arkiv, FTP, etc.)WordWrap	OnClickDDExtLabelClick  TLabelDDExtDisabledLabelLeft#Top� Width:Height6AnchorsakLeftakTopakRight AutoSizeCaption�M�jligg�r nerladdningar till valfri destination (vanliga mappar, ZIP-arkiv, FTP, etc.). Filer laddas f�rst ner till en tempor�r mapp och flyttas d�refter till destinationen.WordWrap	OnClickDDExtLabelClick  TRadioButtonDDExtEnabledButtonLeftTop0WidthLHeightAnchorsakLeftakTopakRight CaptionAnv�nd &skaltill�ggTabOrderOnClickControlChange  TRadioButtonDDExtDisabledButtonLeftTop|WidthDHeightAnchorsakLeftakTopakRight CaptionAnv�nd &tempor�r mappTabOrderOnClickControlChange  TPanelDDExtDisabledPanelLeft"Top� Width;Height3
BevelOuterbvNoneTabOrder
DesignSize;3  	TCheckBoxDDWarnLackOfTempSpaceCheckLeft TopWidth;HeightAnchorsakLeftakTopakRight Caption(&Varna vid otillr�ckligt med diskutrymmeTabOrder OnClickControlChange  	TCheckBoxDDWarnOnMoveCheckLeft TopWidth;HeightAnchorsakLeftakTopakRight Caption%Varna vid &flytt via tempor�r katalogTabOrderOnClickControlChange   	TCheckBoxDDAllowMoveInitCheckLeftTopWidthLHeightAnchorsakLeftakTopakRight Caption<Till�t f&lyttning fr�n fj�rrkatalog till andra applikationerTabOrder OnClickControlChange    	TTabSheet
QueueSheetTagHintBakgrundHelpType	htKeywordHelpKeywordui_pref_backgroundCaptionQue
ImageIndex
TabVisible
DesignSizeua  	TGroupBox
QueueGroupLeftTopWidtheHeight� AnchorsakLeftakTopakRight Caption�verf�ringar i bakgrundenTabOrder  TLabelLabel5LeftTopWidth� HeightCaption'&Maximalt antal samtidiga �verf�ringar:FocusControlQueueTransferLimitEdit  TUpDownEditQueueTransferLimitEditLeftTopWidthIHeight	AlignmenttaRightJustifyMaxValue	MinValueValue	MaxLengthTabOrder   	TCheckBoxQueueAutoPopupCheckLeftTopzWidthQHeightCaptionAVisa bakgrunds�verf�ringarnas prompt &automatiskt vid inaktivitetTabOrder  	TCheckBox
QueueCheckLeftTop2WidthQHeightCaption"&�verf�r som standard i bakgrundenTabOrder  	TCheckBoxRememberPasswordCheckLeftTop� WidthQHeightCaption<Kom ih�g &huvudsessionens l�senord vid bakgrunds�verf�ringarTabOrder  	TCheckBoxQueueNoConfirmationCheckLeftTopbWidthQHeightCaption-I&ngen bekr�ftelser f�r bakgrunds�verf�ringarTabOrder  	TCheckBoxQueueIndividuallyCheckLeftTopJWidthQHeightCaption.&L�gg till varje fil individuellt som standardTabOrder   	TGroupBoxQueueViewGroupLeftTop� WidtheHeightcAnchorsakLeftakTopakRight CaptionK�listaTabOrder TRadioButtonQueueViewShowButtonLeftTopWidthQHeightCaptionVi&saTabOrder   TRadioButtonQueueViewHideWhenEmptyButtonLeftTop-WidthQHeightCaption&D�lj ifall tomTabOrder  TRadioButtonQueueViewHideButtonLeftTopEWidthQHeightCaption&D�ljTabOrder    	TTabSheetStorageSheetTagHintLagringHelpType	htKeywordHelpKeywordui_pref_storageCaptionStor
ImageIndex
TabVisible
DesignSizeua  	TGroupBoxStorageGroupLeftTopWidtheHeightHAnchorsakLeftakTopakRight CaptionInst�llningar f�r lagringTabOrder  TRadioButtonRegistryStorageButtonLeftTopWidth!HeightCaptionWindowsre&gistretTabOrder OnClickControlChange  TRadioButtonIniFileStorageButton2LeftTop-Width!HeightCaption&INI-fil (winscp.ini)TabOrderOnClickControlChange   	TGroupBoxTemporaryDirectoryGrouoLeftTopXWidtheHeight� AnchorsakLeftakTopakRight CaptionTempor�r katalogTabOrder
DesignSizee�   TLabelLabel6LeftTopWidthDHeightAnchorsakLeftakTopakRight AutoSizeCaption>Ange var nerladdade och redigerade filer ska sparas tempor�rt.WordWrap	  TRadioButton DDSystemTemporaryDirectoryButtonLeftTop-Width)HeightCaption#&Anv�nd systemets tempor�ra katalogTabOrder OnClickControlChange  TRadioButton DDCustomTemporaryDirectoryButtonLeftTopEWidth� HeightCaptionAnv�nd den h�r &katalogen:TabOrderOnClickControlChange  TDirectoryEditDDTemporaryDirectoryEditLeft� TopAWidth� HeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPathEditAfterDialog
DialogText.V�lj katalog f�r tempor�ra dra && sl�pp filer.ClickKey@AnchorsakLeftakTopakRight TabOrderTextDDTemporaryDirectoryEditOnClickControlChange  	TCheckBoxTemporaryDirectoryCleanupCheckLeftTop� WidthEHeightAnchorsakLeftakTopakRight Caption-&Rensa gamla tempor�ra kataloger vid uppstartTabOrderOnClickControlChange  	TCheckBox%ConfirmTemporaryDirectoryCleanupCheckLeft Top� Width5HeightAnchorsakLeftakTopakRight Caption&Fr�ga innan rensningTabOrderOnClickControlChange  	TCheckBox$TemporaryDirectoryAppendSessionCheckLeftTop^WidthEHeightAnchorsakLeftakTopakRight Caption/L�gg till &sessionsnamn till tempor�ra s�kv�genTabOrderOnClickControlChange  	TCheckBox!TemporaryDirectoryAppendPathCheckLeftTopwWidthEHeightAnchorsakLeftakTopakRight Caption.L�gg till f&j�rrs�kv�g till tempor�ra s�kv�genTabOrderOnClickControlChange   	TGroupBoxOtherStorageGroupLeftTop%WidtheHeight5AnchorsakLeftakTopakRight Caption�vrigtTabOrder
DesignSizee5  TLabelRandomSeedFileLabelLeftTopWidthUHeightCaptionSl&umpfr�fil:FocusControlRandomSeedFileEdit  TFilenameEditRandomSeedFileEditLeft� TopWidth� HeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPathEditAfterDialog
DefaultExtlogFilter/Slumpfr�filer (*.rnd|*.rnd|Alla filer (*.*)|*.*DialogOptionsofHideReadOnlyofPathMustExist DialogTitleV�lj fil f�r slumpfr�OnCreateEditDialog"RandomSeedFileEditCreateEditDialogClickKey@AnchorsakLeftakTopakRight TabOrder TextRandomSeedFileEditOnChangeControlChange    	TTabSheetTransferEnduranceSheetTagHintToleransHelpType	htKeywordHelpKeywordui_pref_resumeCaptionEndur
ImageIndex
TabVisible
DesignSizeua  	TGroupBox	ResumeBoxLeftTopWidtheHeight{AnchorsakLeftakTopakRight Caption:Aktivera �verf�ringspaus/�verf�r till tempor�r filnamn f�rTabOrder  TLabelResumeThresholdUnitLabelLeft� TopGWidthHeightCaptionKiBFocusControlResumeThresholdEdit  TRadioButtonResumeOnButtonLeftTopWidthIHeightCaptionA&lla filerTabOrder OnClickControlChange  TRadioButtonResumeSmartButtonLeftTop-Width� HeightCaptionFiler st�&rre �n:TabOrderOnClickControlChange  TRadioButtonResumeOffButtonLeftTop]WidthIHeightCaptionA&vaktiveraTabOrderOnClickControlChange  TUpDownEditResumeThresholdEditLeft-TopCWidthTHeight	AlignmenttaRightJustify	Increment
MaxValue  @ TabOrderOnClickControlChange   	TGroupBoxSessionReopenGroupLeftTop� WidtheHeight� AnchorsakLeftakTopakRight CaptionAutomatisk �teranslutningTabOrder TLabelSessionReopenAutoLabelLeft"TopHWidthPHeightCaption&�teranslut efter:FocusControlSessionReopenAutoEdit  TLabelSessionReopenAutoSecLabelLeft� TopHWidth(HeightCaptionsekunderFocusControlSessionReopenAutoEdit  TLabelSessionReopenTimeoutLabelLeft"TopdWidthlHeightCaption&Forts�tt �teransluta i:FocusControlSessionReopenTimeoutEdit  TLabelSessionReopenTimeoutSecLabelLeft� TopdWidth(HeightCaptionsekunderFocusControlSessionReopenTimeoutEdit  	TCheckBoxSessionReopenAutoCheckLeftTopWidthQHeightCaption>&Automatiskt �teranslut session, om den bryts under �verf�ringTabOrder OnClickControlChange  TUpDownEditSessionReopenAutoEditLeft� TopCWidthQHeight	AlignmenttaRightJustify	IncrementMaxValue,MinValueValue	MaxLengthTabOrder  	TCheckBoxSessionReopenAutoIdleCheckLeftTop-WidthQHeightCaption8&Automatiskt �teranslut session, om den bryts under idleTabOrderOnClickControlChange  TUpDownEditSessionReopenTimeoutEditLeft� Top_WidthQHeight	AlignmenttaRightJustify	IncrementMaxValue�Q 	MaxLengthTabOrder
OnGetValue SessionReopenTimeoutEditGetValue
OnSetValue SessionReopenTimeoutEditSetValue    	TTabSheetUpdatesSheetTagHintUppdateringarHelpType	htKeywordHelpKeywordui_pref_updatesCaptionUpd
ImageIndex
TabVisible
DesignSizeua  	TGroupBoxUpdatesGroupLeftTopWidtheHeight{AnchorsakLeftakTopakRight Caption1Kontrollera automatisk om det finns uppdateringarTabOrder  TRadioButtonUpdatesNeverButtonLeftTopWidthIHeightCaptionAldrigTabOrder OnClickControlChange  TRadioButtonUpdatesDailyButtonLeftTop-Width� HeightCaptionDagligenTabOrderOnClickControlChange  TRadioButtonUpdatesWeeklyButtonLeftTopEWidth� HeightCaptionVeckovisTabOrderOnClickControlChange  TRadioButtonUpdatesMonthlyButtonLeftTop]Width� HeightCaption	M�nadsvisTabOrderOnClickControlChange   	TGroupBoxUpdatesProxyGroupLeftTop� WidtheHeight� AnchorsakLeftakTopakRight Caption
AnslutningTabOrder
DesignSizee�   TLabelUpdatesProxyHostLabelLeft"Top[WidthQHeightCaptionProxy &v�rdnamn:FocusControlUpdatesProxyHostEdit  TLabelUpdatesProxyPortLabelLeft� Top[Width<HeightAnchorsakTopakRight CaptionPo&rtnummer:FocusControlUpdatesProxyPortEdit  TUpDownEditUpdatesProxyPortEditLeft� ToplWidth^Height	AlignmenttaRightJustifyMaxValue��  MinValueValueAnchorsakTopakRight TabOrder  TEditUpdatesProxyHostEditLeft"ToplWidth� HeightAnchorsakLeftakTopakRight 	MaxLength2TabOrderTextUpdatesProxyHostEdit  TRadioButtonUpdatesProxyCheckLeftTopEWidthMHeightCaptionA&nv�nd proxyserverTabOrderOnClickControlChange  TRadioButtonUpdatesDirectCheckLeftTopWidthMHeightCaptionIngen &proxyTabOrder OnClickControlChange  TRadioButtonUpdatesAutoCheckLeftTop-WidthMHeightCaption(Detektera &automatisk proxyinst�llningarTabOrderOnClickControlChange   	TGroupBoxUpdatesOptionsGroupLeftTop� WidtheHeight3AnchorsakLeftakTopakRight Caption
AlternativTabOrder
DesignSizee3  TLabelLabel10LeftTopWidthsHeightCaption+Kontrollera ifall det finns &betaversioner:FocusControlUpdatesBetaVersionsCombo  	TComboBoxUpdatesBetaVersionsComboLeftTopWidth=HeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeightTabOrder     	TTabSheetCopyParamListSheetTagHintF�rinst�llningarHelpType	htKeywordHelpKeywordui_pref_presetsCaptionPres
ImageIndex
TabVisible
DesignSizeua  	TGroupBoxCopyParamListGroupLeftTopWidtheHeightAnchorsakLeftakTopakRight Caption�verf�r f�rinst�llningarTabOrder 
DesignSizee  	TListViewCopyParamListViewLeftTopWidthDHeight� AnchorsakLeftakTopakRightakBottom ColumnsCaptionBeskrivning f�rinst�llningarWidthd Caption
AutomatiskTagWidth(  ColumnClickDragModedmAutomaticHideSelection	OwnerData	ReadOnly		RowSelect	ParentShowHintShowHint	TabOrder 	ViewStylevsReportOnDataCopyParamListViewData
OnDblClickCopyParamListViewDblClick	OnEndDragListViewEndDrag
OnDragDropCopyParamListViewDragDrop
OnDragOverListViewDragOver	OnInfoTipCopyParamListViewInfoTip	OnKeyDownCopyParamListViewKeyDownOnSelectItemListViewSelectItemOnStartDragListViewStartDrag  TButtonAddCopyParamButtonLeftTop� WidthSHeightAnchorsakRightakBottom Caption&L�gg till...TabOrderOnClickAddEditCopyParamButtonClick  TButtonRemoveCopyParamButtonLeftTop� WidthSHeightAnchorsakRightakBottom Caption&Ta bortTabOrderOnClickRemoveCopyParamButtonClick  TButtonUpCopyParamButtonLeftTop� WidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickUpDownCopyParamButtonClick  TButtonDownCopyParamButtonLeftTop� WidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickUpDownCopyParamButtonClick  TButtonEditCopyParamButtonLeftpTop� WidthSHeightAnchorsakRightakBottom Caption&Redigera...TabOrderOnClickAddEditCopyParamButtonClick  TButtonDuplicateCopyParamButtonLeftpTop� WidthSHeightAnchorsakRightakBottom Caption&Dubblera...TabOrderOnClickAddEditCopyParamButtonClick   	TGroupBoxCopyParamListOptionsGroupLeftTop$WidtheHeight3AnchorsakLeftakTopakRightakBottom Caption
AlternativTabOrder 	TCheckBoxCopyParamAutoSelectNoticeCheckLeftTopWidthQHeightCaptionQ&Visa meddelanden n�r f�rinst�llda �verf�ringsinst�llningar har valts automatisktTabOrder OnClickControlChange    	TTabSheetWindowSheetTagHintF�nsterHelpType	htKeywordHelpKeywordui_pref_windowCaptionWin
ImageIndex
TabVisible
DesignSizeua  	TGroupBoxPathInCaptionGroupLeftTopWidtheHeight^AnchorsakLeftakTopakRight CaptionS�kv�g i f�nstertitelTabOrder  TRadioButtonPathInCaptionFullButtonLeftTopWidthQHeightCaptionVisa &l�ng s�kv�gTabOrder   TRadioButtonPathInCaptionShortButtonLeftTop,WidthQHeightCaptionVisa &kort s�kv�gTabOrder  TRadioButtonPathInCaptionNoneButtonLeftTopCWidthQHeightCaption
Visa &inteTabOrder   	TGroupBoxWindowMiscellaneousGroupLeftToplWidtheHeight5AnchorsakLeftakTopakRight Caption�vrigtTabOrder
DesignSizee5  	TCheckBoxMinimizeToTrayCheckLeftTopWidthEHeightAnchorsakLeftakTopakRight CaptionJ&Minimera huvudf�nstret till aktivitetsf�ltets statusomr�de (systemf�ltet)TabOrder OnClickControlChange    	TTabSheetSecuritySheetTagHintS�kerhetHelpType	htKeywordHelpKeywordui_pref_securityCaptionSecurity
ImageIndex
TabVisible
DesignSizeua  	TGroupBoxMasterPasswordGroupLeftTopWidtheHeight\AnchorsakLeftakTopakRight CaptionHuvudl�senordTabOrder 
DesignSizee\  TButtonSetMasterPasswordButtonLeftTop3WidthEHeightAnchorsakLeftakTopakRight Caption�&ndra huvudl�senord...TabOrderOnClickSetMasterPasswordButtonClick  	TCheckBoxUseMasterPasswordCheckLeftTopWidthKHeightAnchorsakLeftakTopakRight CaptionAn&v�nd huvudl�senordTabOrder OnClickUseMasterPasswordCheckClick    	TTabSheetIntegrationAppSheetTagHintApplikationerHelpType	htKeywordHelpKeywordui_pref_integration_appCaptionIntgApp
ImageIndex
TabVisible
DesignSizeua  	TGroupBoxExternalAppsGroupLeftTopWidtheHeight� AnchorsakLeftakTopakRight CaptionExterna applikationerTabOrder 
DesignSizee�   TLabelLabel2LeftTopWidth=HeightCaptionS�kv�g till &PuTTY:FocusControlPuttyPathEdit  TEditPuttyPathEditLeftTop&WidthJHeightAnchorsakLeftakTopakRight TabOrder TextPuttyPathEditOnChangeControlChange  	TCheckBoxPuttyPasswordCheck2LeftTopaWidthAHeightCaption;&Kom ih�g sessionsl�senord och �verf�r det till PuTTY (SSH)TabOrder  	TCheckBoxAutoOpenInPuttyCheckLeftTop� WidthAHeightCaption(&�ppna automatiskt en ny session i PuTTYTabOrder  TButtonPuttyPathBrowseButtonLeft� TopAWidthKHeightAnchorsakTopakRight Caption&Bl�ddra...TabOrderOnClickPuttyPathBrowseButtonClick  TButtonPuttyPathResetButtonLeftTopAWidthAHeightAnchorsakTopakRight Caption
�t&erst�llTabOrderOnClickPuttyPathResetButtonClick  	TCheckBoxTelnetForFtpInPuttyCheckLeftTopzWidthAHeightCaption0�ppna &Telnetsessioner i PuTTY f�r FTP-sessionerTabOrder     TPanel	LeftPanelLeft Top Width� HeightkAlignalLeft
BevelOuterbvNoneTabOrder 
DesignSize� k  	TTreeViewNavigationTreeLeftTop	WidthtHeightaAnchorsakLeftakTopakRightakBottom HideSelectionHotTrack	IndentReadOnly	ShowButtonsShowRootTabOrder OnChangeNavigationTreeChangeOnCollapsingNavigationTreeCollapsing
Items.Data
�  	   %          ��������       EnvironmentX#          ��������        
InterfaceX           ��������        WindowX           ��������        PanelsX#          ��������        
CommanderX"          ��������        	ExplorerX           ��������        EditorX"          ��������       	TransferX!          ��������        PresetsX"          ��������        	DragDropX$          ��������        BackgroundX           ��������        ResumeX"          ��������        	SecurityX!          ��������        LoggingX%       	   ��������       IntegrationX&          ��������        ApplicationsX"       
   ��������        	CommandsX!          ��������        StorageX!          ��������        UpdatesX    TButton
HelpButtonLeft�TopqWidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrderOnClickHelpButtonClick  TButtonExportButtonLeftTopqWidthKHeightAnchorsakLeftakBottom CaptionE&xportera...TabOrderOnClickExportButtonClick   TPF0TProgressFormProgressFormLeft�Top#HelpType	htKeywordHelpKeywordui_progressBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption	OperationClientHeight� ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrderPositionpoMainFormCenterOnHideFormHideOnShowFormShow
DesignSize��  PixelsPerInch`
TextHeight TLabelOnceDoneOperationLabelLeftBTopXWidthDHeightCaptionN�r &f�rdig:FocusControlOnceDoneOperationCombo  TAnimateAnimateLeft
TopWidth-Height<ActiveAnchorsakLeftakTopakRight AutoSize	StopFrame  TButtonCancelButtonLeft@TopWidthPHeightAnchorsakTopakRight Cancel	CaptionAvbrytTabOrder OnClickCancelButtonClick  TButtonMinimizeButtonLeft@Top(WidthPHeightAnchorsakTopakRight Caption	&MinimeraTabOrderOnClickMinimizeButtonClick  TPanel	MainPanelLeft
TopAWidth-HeightDAnchorsakLeftakTopakRight 
BevelOuterbvNoneTabOrder
DesignSize-D  TLabelLabel1Left TopWidthHeightCaptionFil:  
TPathLabel	FileLabelLeft8TopWidth� HeightIndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TLabelTargetLabelLeft TopWidth"HeightCaptionM�l:  
TPathLabelTargetPathLabelLeft8TopWidth� HeightIndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TProgressBarTopProgressLeft Top*Width-HeightAnchorsakLeftakTopakRight Min MaxdParentShowHintShowHint	TabOrder    TPanelTransferPanelLeft
Top� Width-Height?AnchorsakLeftakTopakRight 
BevelOuterbvNoneTabOrder
DesignSize-?  TLabelStartTimeLabelLeftXTopWidthAHeight	AlignmenttaRightJustifyAutoSizeCaption00:00:00  TLabelTimeLeftLabelLeftXTopWidthAHeight	AlignmenttaRightJustifyAutoSizeCaption00:00:00  TLabelTimeLeftLabelLabelLeft TopWidth+HeightCaption	Tid kvar:  TLabelCPSLabelLeft� TopWidthAHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption0 KiB/s  TLabelTimeElapsedLabelLeft� TopWidthAHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption00:00:00  TLabelBytesTransferedLabelLeftXTopWidthAHeight	AlignmenttaRightJustifyAutoSizeCaption0 KiB  TLabelLabel3Left� TopWidthBHeightAnchorsakTopakRight CaptionF�rfluten tid:  TLabelStartTimeLabelLabelLeft TopWidth/HeightCaption
Start tid:  TLabelLabel4Left TopWidthRHeightCaptionBytes �verf�rda:  TLabelLabel12Left� TopWidth"HeightAnchorsakTopakRight Caption
Hastighet:  TProgressBarBottomProgressLeft Top%Width-HeightAnchorsakLeftakTopakRight Min MaxdParentShowHintShowHint	TabOrder    TPanel
SpeedPanelLeft:Top� Width\Height)AnchorsakTopakRight 
BevelOuterbvNoneTabOrder TLabelSpeedLabel2LeftTop WidthEHeightCaption&Hastighet (KiB/s)FocusControl
SpeedCombo  THistoryComboBox
SpeedComboLeftTopWidthPHeightAutoComplete
ItemHeightTabOrder Text
SpeedComboOnExitSpeedComboExit
OnKeyPressSpeedComboKeyPressOnSelectSpeedComboSelectItems.Strings	Unlimited10245122561286432168    	TComboBoxOnceDoneOperationComboLeft@TophWidthPHeightAutoCompleteStylecsDropDownList
ItemHeightTabOrder	OnCloseUpOnceDoneOperationComboCloseUpOnSelectOnceDoneOperationComboSelectItems.StringsF�rbli idleKoppla ifr�nSt�ng av dator   TTimerUpdateTimerEnabledOnTimerUpdateTimerTimerLeftPTop�       TPF0TPropertiesDialogPropertiesDialogLeft�Top� HelpType	htKeywordHelpKeywordui_propertiesBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption
PropertiesClientHeight�ClientWidtheColor	clBtnFace
ParentFont	OldCreateOrder	PositionpoMainFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSizee� PixelsPerInch`
TextHeight TButtonOkButtonLeftcTop�WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top�WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TPageControlPageControlLeftTopWidthZHeightv
ActivePageCommonSheetAnchorsakLeftakTopakRightakBottom TabIndex TabOrder OnChangePageControlChange 	TTabSheetCommonSheetCaptionAllm�nt
DesignSizeRZ  TImageFilesIconImageLeftTopWidth Height Picture.Data
�  TBitmapv  BMv      v   (                    �  �          ��� ��� �� ���  Ɓ  �   w  T  N�  �  w                 3           3333""""""""""3333DDDDDDDDDB 333DDDDDDDDDB333DDDDDDDDDB 33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDD  33DDDDDDDBB33DDDDDDD!  33DDDDDDDBB33DDDDDDD!  33DDDDDDDB333!3333DDDDDDD33333333333DDDDDDD33333333333Transparent	  TBevelBevel1LeftTop/Width@Height	AnchorsakLeftakTopakRight Shape	bsTopLine  TLabelLabel1LeftTop:Width,HeightCaptionPlats:  
TPathLabelLocationLabelLeftUTop:Width� HeightUnixPath	IndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TLabel	FileLabelLeftUTopWidth� HeightAutoSizeCaption	FileLabel  TLabelLabel2LeftTopPWidthHeightCaptionStorlek:  TLabel	SizeLabelLeftUTopPWidth� HeightAnchorsakLeftakTopakRight AutoSizeCaption	SizeLabel  TLabelLinksToLabelLabelLeftTopfWidth(HeightCaptionL�nkar till:  
TPathLabelLinksToLabelLeftXTopfWidth� HeightUnixPath	IndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TBevelBevel2LeftTop}Width@Height	AnchorsakLeftakTopakRight Shape	bsTopLine  TLabelLabel3LeftTop� Width:HeightCaptionFilr�ttigheter:FocusControlRightsFrame  TBevelBevel3LeftTop� Width@Height	AnchorsakLeftakTopakRight Shape	bsTopLine  TLabelLabel4LeftTop� Width HeightCaptionGrupp:FocusControlGroupComboBox  TLabelLabel5LeftTop� Width"HeightCaption�gare:FocusControlOwnerComboBox  TImageFileIconImageLeftTopWidth Height   TBevelRecursiveBevelLeftTop8Width@Height	AnchorsakLeftakTopakRight Shape	bsTopLine  �TRightsExtFrameRightsFrameLeftTTop� Width� HeightmTabOrder  	TComboBoxGroupComboBoxLeftUTop� Width� Height
ItemHeight	MaxLength2TabOrderTextGroupComboBoxOnChangeControlChangeOnExitGroupComboBoxExit  	TComboBoxOwnerComboBoxLeftUTop� Width� Height
ItemHeight	MaxLength2TabOrderTextOwnerComboBoxOnChangeControlChangeOnExitOwnerComboBoxExit  	TCheckBoxRecursiveCheckLeftTopBWidth=HeightAnchorsakLeftakTopakRight Caption/S�tt grupp, �gare och filr�ttigheter &rekursivtTabOrderOnClickControlChange  TButtonCalculateSizeButtonLeft� TopHWidthPHeightAnchorsakTopakRight CaptionB&er�knaTabOrder OnClickCalculateSizeButtonClick   	TTabSheetChecksumSheetCaptionKontrollsumma
ImageIndex
DesignSizeRZ  TLabelLabel6LeftTopWidth.HeightCaption
&Algoritm:FocusControlChecksumAlgEdit  	TListViewChecksumViewLeftTop(WidthFHeight)AnchorsakLeftakTopakRightakBottom ColumnsCaptionFilWidth�	WidthType�  CaptionKontrollsummaWidth�	WidthType�   ColumnClickMultiSelect	ReadOnly		RowSelect		PopupMenuListViewMenuTabOrder	ViewStylevsReportOnContextPopupChecksumViewContextPopup  	TComboBoxChecksumAlgEditLeftPTop	WidthyHeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeight	MaxLength� TabOrder OnChangeChecksumAlgEditChangeItems.Stringsmd5sha1sha224sha256sha384sha512crc32   TButtonChecksumButtonLeft� TopWidthzHeightAnchorsakTopakRight CaptionB&er�kna kontrollsummaTabOrderOnClickChecksumButtonClick  	TGroupBoxChecksumGroupLeftTop(WidthFHeight)AnchorsakLeftakRightakBottom CaptionKontrollsummaTabOrder
DesignSizeF)  TEditChecksumEditLeft
TopWidth2HeightTabStopAnchorsakLeftakTopakRight BorderStylebsNoneColor	clBtnFaceReadOnly	TabOrder TextChecksumEdit     TButton
HelpButtonLeftTop�WidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrderOnClickHelpButtonClick  
TPopupMenuListViewMenuLeftTop� 	TMenuItemCopyCaption&KopieraOnClick	CopyClick    TPF0TRemoteTransferDialogRemoteTransferDialogLeft(Top� HelpType	htKeywordHelpKeywordtask_move_duplicateBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionRemoteTransferDialogClientHeight� ClientWidthJColor	clBtnFace
ParentFont	OldCreateOrderPositionpoMainFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSizeJ�  PixelsPerInch`
TextHeight 	TGroupBoxSymlinkGroupLeftTopWidth:Height� AnchorsakLeftakTopakRightakBottom TabOrder 
DesignSize:�   TLabelSessionLabelLeftTopWidthHHeightCaptionM�l&session:FocusControlSessionCombo  TLabelLabel2LeftTop@WidthpHeightCaptionM�l f�r fj�rr&katalog:FocusControlDirectoryEdit  	TComboBoxSessionComboLeftTop Width$HeightStylecsDropDownListAnchorsakLeftakTopakRight 
ItemHeight	MaxLength� TabOrder OnChangeSessionComboChange  THistoryComboBoxDirectoryEditLeftTopPWidth$HeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeight	MaxLength� TabOrderOnChangeControlChange  	TCheckBoxNotDirectCopyCheckLeftTopmWidth HeightAnchorsakLeftakTopakRight Caption!Dubblera via lokal tempor�r kopiaTabOrderOnClickNotDirectCopyCheckClick   TButtonOkButtonLeftNTop� WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top� WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeft� Top� WidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrderOnClickHelpButtonClick    TPF0�TRightsExtFrameRightsExtFrameWidth� Heightm �TLabel
OctalLabelLeftTopDWidthHeightCaptionO&ktal:FocusControl	OctalEdit  �TGrayedCheckBoxGroupReadCheckTabOrder  �TGrayedCheckBoxGroupWriteCheckTabOrder  �TGrayedCheckBoxGroupExecuteCheckTabOrder  �TGrayedCheckBoxOthersReadCheckTabOrder  �TGrayedCheckBoxOthersWriteCheckTabOrder	  �TGrayedCheckBoxOthersExecuteCheckTabOrder
  �	TCheckBoxDirectoriesXCheckTopYTabOrder  �TEdit	OctalEditLeft7Top@Width@Height	MaxLengthTabOrderText	OctalEditOnChangeOctalEditChangeOnExitOctalEditExit  �TGrayedCheckBoxSetUidCheckTag Left� TopWidthFHeightCaptionS�tt UIDTabOrderOnClickControlChange  �TGrayedCheckBoxSetGIDCheckTag Left� TopWidthFHeightCaptionS�tt GIDTabOrderOnClickControlChange  �TGrayedCheckBoxStickyBitCheckTag Left� Top+WidthFHeightCaption
Sticky bitTabOrderOnClickControlChange  �TButtonCloseButtonLeft� TopPWidthKHeightCaptionSt�ngTabOrderVisibleOnClickCloseButtonClick   TPF0TRightsFrameRightsFrameLeft Top Width� HeightWTabOrder OnContextPopupFrameContextPopup TLabel
OwnerLabelLeftTopWidthHeightCaption&�gareFocusControlOwnerReadCheck  TLabel
GroupLabelLeftTopWidthHeightCaption&GruppFocusControlGroupReadCheck  TLabelOthersLabelLeftTop,WidthHeightCaptionA&ndraFocusControlOthersReadCheck  TSpeedButtonOthersButtonTagLeft Top)Width8HeightFlat	OnClickRightsButtonsClick  TSpeedButtonGroupButtonTagLeft TopWidth8HeightFlat	OnClickRightsButtonsClick  TSpeedButtonOwnerButtonTagLeft TopWidth8HeightFlat	OnClickRightsButtonsClick  TGrayedCheckBoxOwnerReadCheckTag Left:TopWidth"HeightHintL�sCaptionRParentShowHintShowHint	TabOrder OnClickControlChange  TGrayedCheckBoxOwnerWriteCheckTag� Left_TopWidth"HeightHintSkrivCaptionWParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxOwnerExecuteCheckTag@Left� TopWidthHeightHint	K�r/�ppnaCaptionXParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxGroupReadCheckTag Left:TopWidth"HeightCaptionRParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxGroupWriteCheckTagLeft_TopWidth!HeightCaptionWParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxGroupExecuteCheckTagLeft� TopWidthHeightCaptionXParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxOthersReadCheckTagLeft:Top+Width"HeightCaptionRParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxOthersWriteCheckTagLeft_Top+Width!HeightCaptionWParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxOthersExecuteCheckTagLeft� Top+WidthHeightCaptionXParentShowHintShowHint	TabOrderOnClickControlChange  	TCheckBoxDirectoriesXCheckLeftTopAWidth� HeightCaptionAddera &X till katalogerTabOrder	OnClickControlChange  
TPopupMenuRightsPopupImagesRightsImagesOnPopupRightsPopupPopupLeft� Top; 	TMenuItem	Norights1ActionNoRightsAction  	TMenuItemDefaultrights1ActionDefaultRightsAction  	TMenuItem
Allrights1ActionAllRightsAction  	TMenuItem
Leaveasis1ActionLeaveRightsAsIsAction  	TMenuItemN1Caption-  	TMenuItemCopyAsText1ActionCopyTextAction  	TMenuItemCopyAsOctal1ActionCopyOctalAction  	TMenuItemPaste1ActionPasteAction   TActionListRightsActionsImagesRightsImages	OnExecuteRightsActionsExecuteOnUpdateRightsActionsUpdateLeft� Top TActionNoRightsActionCaptionI&nga r�ttigheter
ImageIndex ShortCutN@  TActionDefaultRightsActionCaptionStan&dardr�ttigheter
ImageIndexShortCutD@  TActionAllRightsActionCaption&Alla r�ttigheter
ImageIndexShortCutA@  TActionLeaveRightsAsIsActionCaption&L�mna of�r�ndradShortCutL@  TActionCopyTextActionCaption&Kopiera som text
ImageIndexShortCutC@  TActionCopyOctalActionCaptionKopiera som &oktalt
ImageIndexShortCutO@  TActionPasteActionCaptionKl&istra in
ImageIndexShortCutV@   
TImageListRightsImagesLeft� Bitmap
&2  IL 	    �������������BM6       6   (   @   0           0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �   �   �   �   �   �   �   �   �   �                                                                                                                                                               �   �   �   �   �   �   �   �   �                           �   ��� ��� ��� ��� ��� ��� ��� ��� �                                                                                                                                                               �   ��� ��� ��� ��� ��� ��� ��� �       ���  �� ���  �� ��� �   ���                         ��� �                                                                                                                                                               �   ��� ���     ��� ���     ��� �        �� ���  �� ���  �� �   ��� ��� ��� ��� ��� ��� ��� ��� �                                                                                                                                                               �   ���         ��� ���     ��� �       ���  �� ���  �� ��� �   ���             ��� �   �   �   �                                                                                                                                           ��� ��� ��� ��� ��� �   ��� ���     ���         ��� �        �� ���  �� ���  �� �   ��� ��� ��� ��� ��� �   ��� �                                                                                                                                               ��� ���     ��� ��� �   ���         ��� ���     ��� �       ���  �� ���  �� ��� �   ��� ��� ��� ��� ��� �   �                                                                                                                                                   ���         ��� ��� �   ��� ��� ��� ��� �   �   �   �        �� ���  �� ���  �� �   �   �   �   �   �   �                                                                                                                                                       ��� ���     ��� ��� �   ��� ��� ��� ��� �   ��� �           ���  �� ���  �� ���  �� ���  �� ���  �� ���  ��                                                                                                                                                     ���         ��� ��� �   ��� ��� ��� ��� �   �                �� ���                                 ��� ���                                                                                                                                                     ��� ��� ��� ���     �   �   �   �   �   �                   ��� ���                                 ���  ��                                                                                                                                                     ��� ��� ��� ���     ���                                      �� ���  ��      ��          ��     ���  �� ���                                                                                                                                                     ��� ��� ��� ���                                                                  ��  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             {{  {{  {{  91!     ZZ {{      91!                             {{  {{  {{  ))     ZZ {{      9)J                     ss9 ss9 ss9 JJ9     JJ9 ss9     ))) kk     kk     kk                                                                             ��  ��  ��  {{  ��  {{  ��  {{  {{  !{�       � ���             ��  ��  ��  {{  ��  {{  ��  {{  {{  !{�                 ��  ��  ��  ss9 ��  ss9 ��  ss9 ss9 s{ s{ s{ kk kk kk                                                                             ZZ   � ��� ��  ��  ZZ BBB 91! {{                              ZZ ��  {{  ��  ��  ZZ BBB )) {{                      JJ9 ��  ss9 ��  ��  ss9 JJ9 JJ9 ss9 �� �� s�� JJ9                                         �   �   �   �   �   �   �   �   �             �   �   � ��� ZZ ��� ��� BBB ZZZ       � ���                         ZZ ��  ZZ ��� ��� BBB cZc                             JJ9 ��  ss9 ss9 ��� JJ9 JJ9 �� s�� ��� JJ9                                         �   ��� ��� ��� ��� ��� ��� ��� �             �   �   � ��� ��� kkk BBB     91!   � ���                             )) )) ��� cZc BBB     ))                             ))) ))) ss9 ss9 JJ9     ))) �� ��� ��� ��� ss9 )))                                 �   ���                     ��� �                 �   �   � ��� ��� ��� ���   �   � ���                                 )) cZc ��� ��� ��� ��� BBB                             ))) JJ9 ��� ��� ��� ��� ))) ��� ��� ��� ��� ss9                                 �   ��� ��� ��� ��� ��� ��� ��� �                     �   �   � ��� ���   �   � ���                                         BBB ��� ��� ��� cZc BBB                                 JJ9 ��� ss9 ��� JJ9 JJ9 ��� ��� ��� ��� )))             ��� ��� ��� ��� ��� �   ���                     ��� �                         �   �   �   �   � ��� BBB                                         cZc ��� ��� ��� ��� BBB                                 JJ9 ��� ��� ��� ��� ))) ��� ��� ��� s�� ���             ���                 �   ��� ��� ��� ��� ��� ��� ��� �                       BBB   �   �   � ��� ��� BBB kkk                                 BBB ��� ��� ��� ��� ��� BBB kkk                         JJ9 ��� ��� ss9 ��� ��� ))) ss9 ��� �{{ ��� JJ9             ��� ��� ��� ��� ��� �   ���         ��� �   �   �   �                         �   �   �   �   � ��� BBB                                         BBB ��� ��� )) ��� BBB                                 ))) ��� ���     ��� ))) ��� ��� ��� ���                 ���                 �   ��� ��� ��� ��� �   ��� �                         �   �   � ��� ���   � ���                                                 BBB ��� cZc                                             JJ9 ��� JJ9     s�� s{ ��� s�� ��� JJ9             ��� ��� ��� ��� ��� �   ��� ��� ��� ��� �   �                     �   �   �   � ��� BBB ��� ���   �   � ���                                         BBB ��� ��� ))                                         ))) ��� ��� ))) s�� �� �� �� �� ��             ���         ���     �   �   �   �   �   �                     �   �   �   � ���                       �   � ���                                                                                                             s�� c�� �� �� �� )))             ��� ��� ��� ���     ���                                       �   � ���                              99   �   � ���                                                  99                                                     ))) s{ s{ s{                     ��� ��� ��� ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         BM>       >   (   @   0         �                      ���                                                                                                                                 ����    ���     � �     �       �       �       �      �      �      �     �     ��    �     ���    ���    ����    ������	�  ���� � ���� ���� ���� ���� ��  � �� � �� ���  ���  ��� �������������������                            TPF0�TScpCommanderFormScpCommanderFormLeft� Top WidthMHeight�HelpType	htKeywordHelpKeywordui_commanderCaptionScpCommanderFormOldCreateOrder	PixelsPerInch`
TextHeight � 	TSplitterSplitterLeft9Top� WidthHeightCursorcrHSplitHinte|Dra f�r att �ndra proportioner p� filpaneler. Dubbelklicka f�r att bredden p� filpanelerna ska lika.ResizeStylersUpdateOnCanResizeSplitterCanResizeOnMovedSplitterMoved  �	TSplitterQueueSplitterTopWidth=  �TTBXDockTopDockWidth=Height�  TTBXToolbarMenuToolbarLeft Top CaptionMenyCloseButtonImagesGlyphsModule.ExplorerImagesMenuBar	
ShrinkModetbsmWrapStretch	TabOrder TTBXSubmenuItemLocalMenuButtonCaption&LokalHelpKeywordui_commander_menu#localHint@�ndra layout f�r lokal panel eller �ndra katalog/enhet som visas TTBXItemTBXItem1Action)NonVisualDataModule.LocalChangePathAction  TTBXSeparatorItemTBXSeparatorItem1HintE  TTBXSubmenuItemTBXSubmenuItem2Caption&G� tillHelpKeywordtask_navigateHintG� till katalog TTBXItemTBXItem2Action&NonVisualDataModule.LocalOpenDirAction  TTBXItemTBXItem3Action/NonVisualDataModule.LocalExploreDirectoryAction  TTBXSeparatorItemTBXSeparatorItem2HintE  TTBXItemTBXItem4Action(NonVisualDataModule.LocalParentDirAction  TTBXItemTBXItem5Action&NonVisualDataModule.LocalRootDirAction  TTBXItemTBXItem6Action&NonVisualDataModule.LocalHomeDirAction  TTBXSeparatorItemTBXSeparatorItem3HintE  TTBXItemTBXItem7Action#NonVisualDataModule.LocalBackAction  TTBXItemTBXItem8Action&NonVisualDataModule.LocalForwardAction   TTBXItemTBXItem9Action&NonVisualDataModule.LocalRefreshAction  TTBXItem	TBXItem10Action*NonVisualDataModule.LocalAddBookmarkAction  TTBXItem	TBXItem11Action.NonVisualDataModule.LocalPathToClipboardAction  TTBXSeparatorItemTBXSeparatorItem4HintE  TTBXSubmenuItemTBXSubmenuItem3Caption&SorteraHelpKeywordui_file_panel#sorting_filesHint�ndra filordning i lokal panel TTBXItem	TBXItem12Action,NonVisualDataModule.LocalSortAscendingAction  TTBXSeparatorItemTBXSeparatorItem5HintE  TTBXItem	TBXItem13Action)NonVisualDataModule.LocalSortByNameAction
GroupIndex	RadioItem	  TTBXItem	TBXItem14Action(NonVisualDataModule.LocalSortByExtAction
GroupIndex	RadioItem	  TTBXItem	TBXItem15Action)NonVisualDataModule.LocalSortByTypeAction
GroupIndex	RadioItem	  TTBXItem	TBXItem16Action,NonVisualDataModule.LocalSortByChangedAction
GroupIndex	RadioItem	  TTBXItem	TBXItem17Action)NonVisualDataModule.LocalSortBySizeAction
GroupIndex	RadioItem	  TTBXItem	TBXItem18Action)NonVisualDataModule.LocalSortByAttrAction
GroupIndex	RadioItem	   TTBXSubmenuItemTBXSubmenuItem4Caption&Visa kolumnerHelpKeywordui_file_panel#selecting_columnsHint#V�lj kolumner som ska visas i panel TTBXItem	TBXItem19Action1NonVisualDataModule.ShowHideLocalNameColumnAction  TTBXItem	TBXItem20Action1NonVisualDataModule.ShowHideLocalSizeColumnAction  TTBXItem	TBXItem21Action1NonVisualDataModule.ShowHideLocalTypeColumnAction  TTBXItem	TBXItem22Action4NonVisualDataModule.ShowHideLocalChangedColumnAction  TTBXItem	TBXItem23Action1NonVisualDataModule.ShowHideLocalAttrColumnAction   TTBXItem
TBXItem221Action%NonVisualDataModule.LocalFilterAction   TTBXSubmenuItemTBXSubmenuItem18Caption&MarkeraHelpKeywordui_commander_menu#markHintKommandon f�r markera TTBXItem
TBXItem107Action#NonVisualDataModule.SelectOneAction  TTBXItem
TBXItem108Action NonVisualDataModule.SelectAction  TTBXItem
TBXItem109Action"NonVisualDataModule.UnselectAction  TTBXItem
TBXItem110Action#NonVisualDataModule.SelectAllAction  TTBXItem
TBXItem111Action)NonVisualDataModule.InvertSelectionAction  TTBXItem
TBXItem112Action(NonVisualDataModule.ClearSelectionAction  TTBXItem	TBXItem27Action*NonVisualDataModule.RestoreSelectionAction   TTBXSubmenuItemTBXSubmenuItem5Caption&FilerHelpKeywordui_commander_menu#filesHintKommandon f�r filoperationer TTBXSubmenuItemTBXSubmenuItem26Caption&NyHelpKeyword
task_indexHintSkapa objekt|Skapa nytt objekt TTBXItem	TBXItem28Action!NonVisualDataModule.NewFileAction  TTBXItem	TBXItem24Action NonVisualDataModule.NewDirAction  TTBXItem
TBXItem209Action!NonVisualDataModule.NewLinkAction   TTBXSeparatorItemTBXSeparatorItem6HintE  TTBXItem	TBXItem25Action%NonVisualDataModule.CurrentOpenAction  TTBXItem	TBXItem26Action%NonVisualDataModule.CurrentEditAction  TTBXSubmenuItemTBXSubmenuItem25Action0NonVisualDataModule.CurrentEditAlternativeAction  TTBXItem	TBXItem29Action%NonVisualDataModule.AddEditLinkAction  TTBXSeparatorItemTBXSeparatorItem7HintE  TTBXItem	TBXItem30Action%NonVisualDataModule.CurrentCopyAction  TTBXItem	TBXItem31Action&NonVisualDataModule.RemoteCopyToAction  TTBXItem	TBXItem32Action%NonVisualDataModule.CurrentMoveAction  TTBXItem	TBXItem33Action&NonVisualDataModule.RemoteMoveToAction  TTBXItem	TBXItem34Action'NonVisualDataModule.CurrentDeleteAction  TTBXItem	TBXItem35Action'NonVisualDataModule.CurrentRenameAction  TTBXItem	TBXItem36ActionNonVisualDataModule.PasteAction  TTBXSeparatorItemTBXSeparatorItem8HintE  TTBXSubmenuItemCustomCommandsMenuAction(NonVisualDataModule.CustomCommandsAction  TTBXSubmenuItemTBXSubmenuItem6Caption&FilnamnHelpKeyword	filenamesHint'Operationer med namn p� vald(a) fil(er) TTBXItem	TBXItem37Action/NonVisualDataModule.FileListToCommandLineAction  TTBXItem	TBXItem38Action-NonVisualDataModule.FileListToClipboardAction  TTBXItem	TBXItem39Action1NonVisualDataModule.FullFileListToClipboardAction  TTBXItem	TBXItem40Action(NonVisualDataModule.UrlToClipboardAction   TTBXSeparatorItemTBXSeparatorItem9HintE  TTBXItem	TBXItem41Action+NonVisualDataModule.CurrentPropertiesAction   TTBXSubmenuItemTBXSubmenuItem7Caption
&KommandonHelpKeywordui_commander_menu#commandsHintAndra kommandon TTBXItem	TBXItem42Action,NonVisualDataModule.CompareDirectoriesAction  TTBXItem	TBXItem43Action%NonVisualDataModule.SynchronizeAction  TTBXItem	TBXItem44Action)NonVisualDataModule.FullSynchronizeAction  TTBXItem	TBXItem45Action-NonVisualDataModule.SynchronizeBrowsingAction  TTBXItem
TBXItem210Action#NonVisualDataModule.FindFilesAction  TTBXSubmenuItemQueueSubmenuItemCaptionK&�HelpKeywordui_queue#managing_the_queueHintKommandon f�r k�listaOnPopupQueueSubmenuItemPopup TTBXItem	TBXItem46Action#NonVisualDataModule.QueueGoToAction  TTBXSeparatorItemTBXSeparatorItem10HintE  TTBXItem	TBXItem47Action(NonVisualDataModule.QueueItemQueryAction  TTBXItem	TBXItem48Action(NonVisualDataModule.QueueItemErrorAction  TTBXItem	TBXItem49Action)NonVisualDataModule.QueueItemPromptAction  TTBXSeparatorItemTBXSeparatorItem11HintE  TTBXItem	TBXItem50Action*NonVisualDataModule.QueueItemExecuteAction  TTBXItem
TBXItem196Action(NonVisualDataModule.QueueItemPauseAction  TTBXItem
TBXItem197Action)NonVisualDataModule.QueueItemResumeAction  TTBXItem	TBXItem51Action)NonVisualDataModule.QueueItemDeleteAction  TTBXComboBoxItemQueueSpeedComboBoxItemAction(NonVisualDataModule.QueueItemSpeedAction  TTBXSeparatorItemTBXSeparatorItem12HintE  TTBXItem	TBXItem52Action%NonVisualDataModule.QueueItemUpAction  TTBXItem	TBXItem53Action'NonVisualDataModule.QueueItemDownAction  TTBXSeparatorItemTBXSeparatorItem48HintE  TTBXSubmenuItemTBXSubmenuItem13Caption&AllaHelpKeywordui_queue#managing_the_queueHint$Administrationskommandon f�r k�massa TTBXItem
TBXItem198Action'NonVisualDataModule.QueuePauseAllAction  TTBXItem
TBXItem199Action(NonVisualDataModule.QueueResumeAllAction    TTBXSeparatorItemTBXSeparatorItem13HintE  TTBXItem	TBXItem54Action!NonVisualDataModule.ConsoleAction  TTBXItem	TBXItem55ActionNonVisualDataModule.PuttyAction  TTBXSeparatorItemTBXSeparatorItem14HintE  TTBXItem	TBXItem56Action(NonVisualDataModule.FileSystemInfoAction  TTBXItem	TBXItem57Action%NonVisualDataModule.ClearCachesAction  TTBXSeparatorItemTBXSeparatorItem15HintE  TTBXItem	TBXItem58Action*NonVisualDataModule.CloseApplicationAction   TTBXSubmenuItemTBXSubmenuItem19Caption&SessionHelpKeywordui_commander_menu#sessionHintKommandon f�r session TTBXItem
TBXItem113Action$NonVisualDataModule.NewSessionAction  TTBXItem
TBXItem218Action*NonVisualDataModule.DuplicateSessionAction  TTBXSubmenuItemTBXSubmenuItem20Action'NonVisualDataModule.SavedSessionsAction  TTBXSeparatorItemTBXSeparatorItem29HintE  TTBXSubmenuItemTBXSubmenuItem21Action(NonVisualDataModule.OpenedSessionsAction  TTBXItem
TBXItem114Action,NonVisualDataModule.SaveCurrentSessionAction  TTBXItem
TBXItem115Action&NonVisualDataModule.CloseSessionAction   TTBXSubmenuItemTBXSubmenuItem9Caption&AlternativHelpKeywordui_commander_menu#optionsHint&�ndra layout/inst�llningar f�r program TTBXSubmenuItemTBXSubmenuItem10Caption&Verktygsf�ltHelpKeywordui_toolbarsHintVisa/d�lj verktygsf�lt TTBXItem	TBXItem59Action.NonVisualDataModule.CommanderToolbarBandAction  TTBXItem	TBXItem60Action.NonVisualDataModule.CommanderSessionBandAction  TTBXItem	TBXItem61Action0NonVisualDataModule.CommanderSelectionBandAction  TTBXItem	TBXItem62Action2NonVisualDataModule.CommanderPreferencesBandAction  TTBXItem	TBXItem63Action+NonVisualDataModule.CommanderSortBandAction  TTBXItem	TBXItem64Action/NonVisualDataModule.CommanderCommandsBandAction  TTBXItem
TBXItem186Action.NonVisualDataModule.CommanderUpdatesBandAction  TTBXItem
TBXItem188Action/NonVisualDataModule.CommanderTransferBandAction  TTBXItem
TBXItem214Action5NonVisualDataModule.CommanderUploadDownloadBandAction  TTBXItem
TBXItem215Action5NonVisualDataModule.CommanderCustomCommandsBandAction  TTBXSeparatorItemTBXSeparatorItem47HintE  TTBXItem
TBXItem191Action&NonVisualDataModule.LockToolbarsAction   TTBXSubmenuItemTBXSubmenuItem11Caption&Lokal panelHelpKeywordui_file_panelHint�ndra layout f�r lokal panel TTBXItem	TBXItem65Action3NonVisualDataModule.CommanderLocalHistoryBandAction  TTBXItem	TBXItem66Action6NonVisualDataModule.CommanderLocalNavigationBandAction  TTBXSeparatorItemTBXSeparatorItem16HintE  TTBXItem	TBXItem67Action#NonVisualDataModule.LocalTreeAction  TTBXSeparatorItemTBXSeparatorItem17HintE  TTBXItem	TBXItem68Action(NonVisualDataModule.LocalStatusBarAction   TTBXSubmenuItemTBXSubmenuItem12CaptionF&j�rrpanelHelpKeywordui_file_panelHint�ndra layout f�r fj�rrpanel TTBXItem	TBXItem69Action4NonVisualDataModule.CommanderRemoteHistoryBandAction  TTBXItem	TBXItem70Action7NonVisualDataModule.CommanderRemoteNavigationBandAction  TTBXSeparatorItemTBXSeparatorItem18HintE  TTBXItem	TBXItem71Action$NonVisualDataModule.RemoteTreeAction  TTBXSeparatorItemTBXSeparatorItem19HintE  TTBXItem	TBXItem72Action)NonVisualDataModule.RemoteStatusBarAction   TTBXSeparatorItemTBXSeparatorItem20HintE  TTBXItem	TBXItem73Action*NonVisualDataModule.CommandLinePanelAction  TTBXItem	TBXItem74Action!NonVisualDataModule.ToolBarAction  TTBXItem	TBXItem75Action#NonVisualDataModule.StatusBarAction  TTBXItem	TBXItem76Action!NonVisualDataModule.ViewLogAction  TTBXSubmenuItemTBXSubmenuItem14CaptionK&�HelpKeywordui_queueHintKonfigurera k�lista TTBXItem	TBXItem77Action#NonVisualDataModule.QueueShowAction	RadioItem	  TTBXItem	TBXItem78Action,NonVisualDataModule.QueueHideWhenEmptyAction	RadioItem	  TTBXItem	TBXItem79Action#NonVisualDataModule.QueueHideAction	RadioItem	  TTBXSeparatorItemTBXSeparatorItem21HintE  TTBXItem	TBXItem80Action&NonVisualDataModule.QueueToolbarAction  TTBXSeparatorItemTBXSeparatorItem22HintE  TTBXSubmenuItemTBXSubmenuItem8Action-NonVisualDataModule.QueueCycleOnceEmptyActionDropdownCombo	 TTBXItem
TBXItem222Action,NonVisualDataModule.QueueIdleOnceEmptyAction	RadioItem	  TTBXItem
TBXItem223Action2NonVisualDataModule.QueueDisconnectOnceEmptyAction	RadioItem	  TTBXItem
TBXItem224Action0NonVisualDataModule.QueueShutDownOnceEmptyAction	RadioItem	   TTBXItem	TBXItem81Action*NonVisualDataModule.QueuePreferencesAction   TTBXSeparatorItemTBXSeparatorItem23HintE  TTBXColorItemColorMenuItemAction#NonVisualDataModule.ColorMenuActionColorclNone TTBXItem
TBXItem216Action&NonVisualDataModule.ColorDefaultAction  TTBXSeparatorItemTBXSeparatorItem50Blank	  TTBXColorPaletteSessionColorPalettePaletteOptionstpoCustomImages OnChangeSessionColorPaletteChange  TTBXSeparatorItemTBXSeparatorItem51HintE  TTBXItem
TBXItem217Action#NonVisualDataModule.ColorPickAction   TTBXSeparatorItemTBXSeparatorItem49HintE  TTBXItem	TBXItem82Action%NonVisualDataModule.PreferencesAction   TTBXSubmenuItemRemoteMenuButtonCaptionF&j�rrHelpKeywordui_commander_menu#remoteHint9�ndra layout f�r fj�rrpanel eller �ndra katalog som visas TTBXItem	TBXItem83Action*NonVisualDataModule.RemoteChangePathAction  TTBXSeparatorItemTBXSeparatorItem24HintE  TTBXSubmenuItemTBXSubmenuItem15Caption&G� tillHelpKeywordtask_navigateHintG� till katalog TTBXItem	TBXItem84Action'NonVisualDataModule.RemoteOpenDirAction  TTBXSeparatorItemTBXSeparatorItem25HintE  TTBXItem	TBXItem85Action)NonVisualDataModule.RemoteParentDirAction  TTBXItem	TBXItem86Action'NonVisualDataModule.RemoteRootDirAction  TTBXItem	TBXItem87Action'NonVisualDataModule.RemoteHomeDirAction  TTBXSeparatorItemTBXSeparatorItem26HintE  TTBXItem	TBXItem88Action$NonVisualDataModule.RemoteBackAction  TTBXItem	TBXItem89Action'NonVisualDataModule.RemoteForwardAction   TTBXItem	TBXItem90Action'NonVisualDataModule.RemoteRefreshAction  TTBXItem	TBXItem91Action+NonVisualDataModule.RemoteAddBookmarkAction  TTBXItem	TBXItem92Action/NonVisualDataModule.RemotePathToClipboardAction  TTBXSeparatorItemTBXSeparatorItem27HintE  TTBXSubmenuItemTBXSubmenuItem16Caption&SorteraHelpKeywordui_file_panel#sorting_filesHint�ndra filordning i fj�rrpanel TTBXItem	TBXItem93Action-NonVisualDataModule.RemoteSortAscendingAction  TTBXSeparatorItemTBXSeparatorItem28HintE  TTBXItem	TBXItem94Action*NonVisualDataModule.RemoteSortByNameAction
GroupIndex	RadioItem	  TTBXItem	TBXItem95Action)NonVisualDataModule.RemoteSortByExtAction
GroupIndex	RadioItem	  TTBXItem
TBXItem193Action*NonVisualDataModule.RemoteSortByTypeAction	RadioItem	  TTBXItem	TBXItem96Action-NonVisualDataModule.RemoteSortByChangedAction
GroupIndex	RadioItem	  TTBXItem	TBXItem97Action*NonVisualDataModule.RemoteSortBySizeAction
GroupIndex	RadioItem	  TTBXItem	TBXItem98Action,NonVisualDataModule.RemoteSortByRightsAction
GroupIndex	RadioItem	  TTBXItem	TBXItem99Action+NonVisualDataModule.RemoteSortByOwnerAction
GroupIndex	RadioItem	  TTBXItem
TBXItem100Action+NonVisualDataModule.RemoteSortByGroupAction
GroupIndex	RadioItem	   TTBXSubmenuItemTBXSubmenuItem17Caption&Visa kolumnerHelpKeywordui_file_panel#selecting_columnsHint#V�lj kolumner som ska visas i panel TTBXItem
TBXItem101Action2NonVisualDataModule.ShowHideRemoteNameColumnAction  TTBXItem
TBXItem102Action2NonVisualDataModule.ShowHideRemoteSizeColumnAction  TTBXItem
TBXItem192Action2NonVisualDataModule.ShowHideRemoteTypeColumnAction  TTBXItem
TBXItem103Action5NonVisualDataModule.ShowHideRemoteChangedColumnAction  TTBXItem
TBXItem104Action4NonVisualDataModule.ShowHideRemoteRightsColumnAction  TTBXItem
TBXItem105Action3NonVisualDataModule.ShowHideRemoteOwnerColumnAction  TTBXItem
TBXItem106Action3NonVisualDataModule.ShowHideRemoteGroupColumnAction  TTBXItem
TBXItem179Action8NonVisualDataModule.ShowHideRemoteLinkTargetColumnAction   TTBXItem
TBXItem220Action&NonVisualDataModule.RemoteFilterAction   TTBXSubmenuItemTBXSubmenuItem22Caption&Hj�lpHelpKeywordui_commander_menu#helpHintHj�lp TTBXItem
TBXItem116Action)NonVisualDataModule.TableOfContentsAction  TTBXSeparatorItemTBXSeparatorItem30HintE  TTBXItem
TBXItem117Action"NonVisualDataModule.HomepageAction  TTBXItem
TBXItem118Action#NonVisualDataModule.ForumPageAction  TTBXItem
TBXItem119Action%NonVisualDataModule.HistoryPageAction  TTBXSeparatorItemTBXSeparatorItem31HintE  TTBXItem
TBXItem120Action)NonVisualDataModule.CheckForUpdatesAction  TTBXSeparatorItemTBXSeparatorItem32HintE  TTBXItem
TBXItem121Action$NonVisualDataModule.DonatePageAction  TTBXSeparatorItemTBXSeparatorItem33HintE  TTBXItem
TBXItem122ActionNonVisualDataModule.AboutAction    TTBXToolbarSelectionToolbarLeft TopNCaption	MarkeringDockPos DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem131Action NonVisualDataModule.SelectAction  TTBXItem
TBXItem132Action"NonVisualDataModule.UnselectAction  TTBXSeparatorItemTBXSeparatorItem37  TTBXItem
TBXItem133Action#NonVisualDataModule.SelectAllAction  TTBXItem
TBXItem134Action)NonVisualDataModule.InvertSelectionAction  TTBXItem
TBXItem135Action(NonVisualDataModule.ClearSelectionAction  TTBXItem
TBXItem200Action*NonVisualDataModule.RestoreSelectionAction   TTBXToolbarPreferencesToolbarLeft Top4CaptionInst�llningarDockPos DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem126Action%NonVisualDataModule.PreferencesAction  TTBXSeparatorItemTBXSeparatorItem36  TTBXItem
TBXItem127Action!NonVisualDataModule.ViewLogAction  TTBXSubmenuItemTBXSubmenuItem24Action)NonVisualDataModule.QueueToggleShowActionDropdownCombo	 TTBXItem
TBXItem128Action#NonVisualDataModule.QueueShowAction	RadioItem	  TTBXItem
TBXItem129Action,NonVisualDataModule.QueueHideWhenEmptyAction	RadioItem	  TTBXItem
TBXItem130Action#NonVisualDataModule.QueueHideAction	RadioItem	    TTBXToolbarSessionToolbarLeft TopCaptionSessionDockModedmCannotFloatDockPos DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	Stretch	TabOrder OnResizeToolBarResizeOnGetBaseSizeToolbarGetBaseSize TTBXItem
TBXItem123Action$NonVisualDataModule.NewSessionAction  TTBXItem
TBXItem219Action*NonVisualDataModule.DuplicateSessionAction  TTBXSeparatorItemTBXSeparatorItem34  TTBXComboBoxItemSessionCombo	EditWidthrDropDownList	MaxVisibleItems  TTBXItem
TBXItem124Action&NonVisualDataModule.CloseSessionAction  TTBXSeparatorItemTBXSeparatorItem35  TTBXSubmenuItemTBXSubmenuItem23Action'NonVisualDataModule.SavedSessionsActionOptionstboDropdownArrow   TTBXItem
TBXItem125Action,NonVisualDataModule.SaveCurrentSessionAction   TTBXToolbarCommandToolbarLeft TophCaptionStandardDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem136Action%NonVisualDataModule.CurrentCopyAction  TTBXItem
TBXItem137Action%NonVisualDataModule.CurrentMoveAction  TTBXSeparatorItemTBXSeparatorItem38  TTBXItem
TBXItem138Action%NonVisualDataModule.CurrentEditAction  TTBXItem
TBXItem139Action%NonVisualDataModule.CurrentOpenAction  TTBXItem
TBXItem140Action'NonVisualDataModule.CurrentRenameAction  TTBXItem
TBXItem141Action'NonVisualDataModule.CurrentDeleteAction  TTBXItem
TBXItem142Action+NonVisualDataModule.CurrentPropertiesAction  TTBXSeparatorItemTBXSeparatorItem39  TTBXItem
TBXItem143Action*NonVisualDataModule.CurrentCreateDirAction  TTBXItem
TBXItem144Action%NonVisualDataModule.AddEditLinkAction   TTBXToolbarSortToolbarLeft Top� CaptionSorteraDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem145Action.NonVisualDataModule.CurrentSortAscendingAction  TTBXSeparatorItemTBXSeparatorItem40  TTBXItem
TBXItem146Action+NonVisualDataModule.CurrentSortByNameAction  TTBXItem
TBXItem147Action*NonVisualDataModule.CurrentSortByExtAction  TTBXItem
TBXItem148Action+NonVisualDataModule.CurrentSortByTypeAction  TTBXItem
TBXItem149Action.NonVisualDataModule.CurrentSortByChangedAction  TTBXItem
TBXItem150Action+NonVisualDataModule.CurrentSortBySizeAction  TTBXItem
TBXItem151Action-NonVisualDataModule.CurrentSortByRightsAction  TTBXItem
TBXItem152Action,NonVisualDataModule.CurrentSortByOwnerAction  TTBXItem
TBXItem153Action,NonVisualDataModule.CurrentSortByGroupAction   TTBXToolbarCommandsToolbarLeft Top� Caption	KommandonDockPos DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem154Action,NonVisualDataModule.CompareDirectoriesAction  TTBXItem
TBXItem155Action%NonVisualDataModule.SynchronizeAction  TTBXItem
TBXItem156Action)NonVisualDataModule.FullSynchronizeAction  TTBXSeparatorItemTBXSeparatorItem41  TTBXItem
TBXItem157Action!NonVisualDataModule.ConsoleAction  TTBXItem
TBXItem190ActionNonVisualDataModule.PuttyAction  TTBXSeparatorItemTBXSeparatorItem42  TTBXItem
TBXItem158Action-NonVisualDataModule.SynchronizeBrowsingAction  TTBXItem
TBXItem227Action#NonVisualDataModule.FindFilesAction   TTBXToolbarUpdatesToolbarLeft Top� CaptionUppdateringarDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXSubmenuItemTBXSubmenuItem1Action%NonVisualDataModule.ShowUpdatesActionDropdownCombo	 TTBXItem
TBXItem184Action)NonVisualDataModule.CheckForUpdatesAction  TTBXSeparatorItemTBXSeparatorItem46HintE  TTBXItem
TBXItem180Action"NonVisualDataModule.HomepageAction  TTBXItem
TBXItem187Action&NonVisualDataModule.DownloadPageAction  TTBXItem
TBXItem181Action#NonVisualDataModule.ForumPageAction  TTBXItem
TBXItem182Action%NonVisualDataModule.HistoryPageAction  TTBXItem
TBXItem185Action$NonVisualDataModule.DonatePageAction  TTBXSeparatorItemTBXSeparatorItem45HintE  TTBXItem
TBXItem183Action,NonVisualDataModule.UpdatesPreferencesAction    TTBXToolbarTransferToolbarLeft(Top� Caption�verf�ringsinst�llningarDockModedmCannotFloatDockPos,DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	Stretch	TabOrderOnResizeToolBarResizeOnGetBaseSizeToolbarGetBaseSize TTBXDropDownItemTransferDropDown	EditWidthrHint*V�lj f�rinst�llda �verf�ringsinst�llningarDropDownList	 TTBXStringListTransferListMaxVisibleItemsMinWidth^  TTBXLabelItemTransferLabelMarginShowAccelChar  TTBXSeparatorItemTBXSeparatorItem52  TTBXItem
TBXItem189Action,NonVisualDataModule.PresetsPreferencesActionDisplayModenbdmImageAndText    TTBXToolbarUploadDownloadToolbarLeft� Top� CaptionUppladdning/NerladdningDockPos� DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder	Visible TTBXItem
TBXItem213Action$NonVisualDataModule.RemoteCopyAction  TTBXItem
TBXItem212Action#NonVisualDataModule.LocalCopyAction   TTBXToolbarCustomCommandsToolbarLeft� Top� CaptionEgna kommandonDockPos� DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder
Visible   �TPanelRemotePanelLeft>Top� Width�HeightConstraints.MinHeight� Constraints.MinWidth� TabOrder � 
TPathLabelRemotePathLabelLeft TopOWidth�HeightUnixPath	HotTrack	OnGetStatusRemotePathLabelGetStatusOnPathClickRemotePathLabelPathClickAutoSize
OnDblClickPathLabelDblClick  �	TSplitterRemotePanelSplitterLeft Top� Width�HeightCursorcrVSplitHint`Dra f�r att �ndra storlek p� katalogtr�d. Dubbelklicka f�r att g�r h�jden p� katalogtr�den lika.AlignalTop  �TTBXStatusBarRemoteStatusBarTop� Width�SimplePanel	  �TUnixDirViewRemoteDirViewLeft Top� Width�HeightaConstraints.MinHeightF
NortonLikenlOnOnUpdateStatusBarRemoteDirViewUpdateStatusBar	PathLabelRemotePathLabelAddParentDir	OnDDFileOperationExecuted(RemoteFileControlDDFileOperationExecutedOnPathChangeRemoteDirViewPathChange  �TUnixDriveViewRemoteDriveViewTop^Width�Height-AlignalTopConstraints.MinHeightHideSelectionTabStop  TTBXDockRemoteTopDockLeft Top Width�HeightOFixAlign	 TTBXToolbarRemoteHistoryToolbarLeft TopCaptionFj�rrhistorikDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXSubmenuItemRemoteBackButtonAction$NonVisualDataModule.RemoteBackActionDropdownCombo	  TTBXSubmenuItemRemoteForwardButtonAction'NonVisualDataModule.RemoteForwardActionDropdownCombo	   TTBXToolbarRemoteNavigationToolbarLeft Top5CaptionFj�rrnavigeringDockPos DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem165Action)NonVisualDataModule.RemoteParentDirAction  TTBXItem
TBXItem166Action'NonVisualDataModule.RemoteRootDirAction  TTBXItem
TBXItem167Action'NonVisualDataModule.RemoteHomeDirAction  TTBXItem
TBXItem168Action'NonVisualDataModule.RemoteRefreshAction  TTBXSeparatorItemTBXSeparatorItem44  TTBXItem
TBXItem170Action$NonVisualDataModule.RemoteTreeAction   TTBXToolbarRemotePathToolbarLeft Top CaptionFj�rrs�kv�g
DockableTodpTopdpBottom DockModedmCannotFloatDockPos ImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	Stretch	TabOrder OnResizeToolBarResizeOnGetBaseSizeToolbarGetBaseSize TTBXComboBoxItemRemotePathComboBox	EditWidth� 	ShowImage	DropDownList	MaxVisibleItemsShowListImages	OnAdjustImageIndex"RemotePathComboBoxAdjustImageIndex
OnDrawItemRemotePathComboBoxDrawItemOnItemClickRemotePathComboBoxItemClickOnMeasureWidthRemotePathComboBoxMeasureWidthOnCancelRemotePathComboBoxCancel  TTBXItem
TBXItem169Action'NonVisualDataModule.RemoteOpenDirAction    TTBXDockRemoteBottomDockLeft Top� Width�Height	FixAlign	PositiondpBottom   �TPanel
QueuePanelTopWidth=HeighttTabOrder �	TListView
QueueView2Width=HeightZTabStop  �TTBXDock	QueueDockWidth=   TPanel
LocalPanelLeft Top� Width9HeightAlignalLeft
BevelOuterbvNoneConstraints.MinHeight� Constraints.MinWidth� TabOrder  
TPathLabelLocalPathLabelLeft TopOWidth9HeightHotTrack	OnGetStatusLocalPathLabelGetStatusOnPathClickLocalPathLabelPathClickAutoSize	PopupMenu#NonVisualDataModule.LocalPanelPopup
OnDblClickPathLabelDblClick  	TSplitterLocalPanelSplitterLeft Top� Width9HeightCursorcrVSplitHint`Dra f�r att �ndra storlek p� katalogtr�d. Dubbelklicka f�r att g�r h�jden p� katalogtr�den lika.AlignalTopAutoSnapMinSizeFResizeStylersUpdate  TTBXStatusBarLocalStatusBarLeft Top� Width9HeightPanels ParentShowHintSimplePanel	ShowHint	UseSystemFontOnClickLocalStatusBarClick  TDirViewLocalDirViewLeft Top� Width9HeightaAlignalClientConstraints.MinHeightFFullDrag	HideSelection	PopupMenu%NonVisualDataModule.LocalDirViewPopupTabOrder	ViewStylevsReportOnColumnRightClickDirViewColumnRightClick	OnEditingDirViewEditingOnEnterLocalDirViewEnterDirColProperties.ExtVisible	PathLabelLocalPathLabelOnUpdateStatusBarLocalDirViewUpdateStatusBarOnGetSelectFilterRemoteDirViewGetSelectFilterHeaderImagesGlyphsModule.ArrowImagesAddParentDir	OnLoadedDirViewLoadedOnDDDragEnterLocalFileControlDDDragEnterOnDDDragLeaveFileControlDDDragLeaveOnDDDragOverLocalFileControlDDDragOverOnDDTargetHasDropHandler"LocalDirViewDDTargetHasDropHandlerOnDDFileOperationLocalFileControlDDFileOperationOnDDMenuPopupLocalFileControlDDMenuPopup
OnExecFileLocalDirViewExecFileOnMatchMaskDirViewMatchMaskOnGetOverlayRemoteDirViewGetOverlayConfirmDeleteWatchForChanges	OnFileIconForNameLocalDirViewFileIconForNameOnHistoryChangeDirViewHistoryChangeOnPathChangeLocalDirViewPathChange  TTBXDockLocalTopDockLeft Top Width9HeightOFixAlign	 TTBXToolbarLocalHistoryToolbarLeft TopCaptionLokal historikDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXSubmenuItemLocalBackButtonAction#NonVisualDataModule.LocalBackActionDropdownCombo	  TTBXSubmenuItemLocalForwardButtonAction&NonVisualDataModule.LocalForwardActionDropdownCombo	   TTBXToolbarLocalNavigationToolbarLeft Top5CaptionLokal navigeringDockPos DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem159Action(NonVisualDataModule.LocalParentDirAction  TTBXItem
TBXItem160Action&NonVisualDataModule.LocalRootDirAction  TTBXItem
TBXItem161Action&NonVisualDataModule.LocalHomeDirAction  TTBXItem
TBXItem162Action&NonVisualDataModule.LocalRefreshAction  TTBXSeparatorItemTBXSeparatorItem43  TTBXItem
TBXItem164Action#NonVisualDataModule.LocalTreeAction   TTBXToolbarLocalPathToolbarLeft Top CaptionLokal s�kv�g
DockableTodpTopdpBottom DockModedmCannotFloatDockPos ImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	Stretch	TabOrder OnResizeToolBarResizeOnGetBaseSizeToolbarGetBaseSize TTBXComboBoxItemLocalPathComboBox	EditWidth� 	ShowImage	DropDownList	MaxVisibleItemsShowListImages	OnAdjustImageIndex!LocalPathComboBoxAdjustImageIndexOnItemClickLocalPathComboBoxItemClickOnCancelLocalPathComboBoxCancel  TTBXItem
TBXItem163Action&NonVisualDataModule.LocalOpenDirAction    
TDriveViewLocalDriveViewLeft Top^Width9Height-WatchDirectory	DirViewLocalDirViewOnRefreshDrivesLocalDriveViewRefreshDrivesOnDDDragEnterLocalFileControlDDDragEnterOnDDDragLeaveFileControlDDDragLeaveOnDDDragOverLocalFileControlDDDragOverOnDDFileOperationLocalFileControlDDFileOperationOnDDMenuPopupLocalFileControlDDMenuPopupAlignalTopConstraints.MinHeightHideSelectionIndentParentColorTabOrderTabStopOnEnterLocalDriveViewEnter  TTBXDockLocalBottomDockLeft Top� Width9Height	FixAlign	PositiondpBottom   TTBXDock
BottomDockLeft Top�Width=Height5FixAlign	PositiondpBottom TTBXToolbarToolbarToolbarLeft TopCaption	KommandonDockPos DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHintStretch	TabOrder  TTBXItem
TBXItem171Action'NonVisualDataModule.CurrentRenameActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem172Action%NonVisualDataModule.CurrentEditActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem173Action%NonVisualDataModule.CurrentCopyActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem174Action%NonVisualDataModule.CurrentMoveActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem175Action*NonVisualDataModule.CurrentCreateDirActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem176Action'NonVisualDataModule.CurrentDeleteActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem177Action+NonVisualDataModule.CurrentPropertiesActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem178Action*NonVisualDataModule.CloseApplicationActionDisplayModenbdmImageAndTextStretch	   TTBXToolbarCommandLineToolbarLeft Top CaptionCommandLineToolbarDockModedmCannotFloatStretch	TabOrderVisibleOnResizeToolBarResizeOnGetBaseSizeToolbarGetBaseSize TTBXLabelItemCommandLinePromptLabelCaption
CommandX >Margin  TTBXComboBoxItemCommandLineComboOnBeginEditCommandLineComboBeginEditExtendedAccept	OnPopupCommandLineComboPopup    TTBXStatusBar	StatusBarLeft Top�Width=ImagesGlyphsModule.SessionImagesPanelsSizedStretchPriorityTag TextTruncationtwEndEllipsis 	AlignmenttaCenter
ImageIndexMaxSize#Size#Tag  	AlignmenttaCenterMaxSizeFViewPrioritybSizeFTag TextTruncationtwEndEllipsis 	AlignmenttaCenter
ImageIndex MaxSize#Size#Tag  	AlignmenttaCenterMaxSizePViewPrioritycSizePTag TextTruncationtwEndEllipsis  ParentShowHint	PopupMenu%NonVisualDataModule.CommanderBarPopupShowHint	UseSystemFontOnPanelDblClickStatusBarPanelDblClick     TPF0�TScpExplorerFormScpExplorerFormLeft� Top� Width�HeightHelpType	htKeywordHelpKeywordui_explorerActiveControlRemoteDirViewCaptionScpExplorerFormOldCreateOrder	PixelsPerInch`
TextHeight �	TSplitterQueueSplitterTopPWidth�  �TTBXDockTopDockWidth�Height�  TTBXToolbarMenuToolbarLeft Top CaptionMenyCloseButtonImagesGlyphsModule.ExplorerImagesMenuBar	
ShrinkModetbsmWrapStretch	TabOrder  TTBXSubmenuItemTBXSubmenuItem5Caption&FilHelpKeywordui_explorer_menu#fileHintFiloperationer TTBXSubmenuItemTBXSubmenuItem26Caption&NyHelpKeyword
task_indexHintSkapa objekt|Skapa nytt objekt TTBXItem
TBXItem135Action!NonVisualDataModule.NewFileAction  TTBXItem
TBXItem136Action NonVisualDataModule.NewDirAction  TTBXItem
TBXItem209Action!NonVisualDataModule.NewLinkAction   TTBXSeparatorItemTBXSeparatorItem20HintE  TTBXItem	TBXItem25Action%NonVisualDataModule.CurrentOpenAction  TTBXItem	TBXItem26Action%NonVisualDataModule.CurrentEditAction  TTBXSubmenuItemTBXSubmenuItem9Action0NonVisualDataModule.CurrentEditAlternativeAction  TTBXItemTBXItem4Action%NonVisualDataModule.AddEditLinkAction  TTBXSeparatorItemTBXSeparatorItem7HintE  TTBXItem	TBXItem34Action'NonVisualDataModule.CurrentDeleteAction  TTBXItem	TBXItem35Action'NonVisualDataModule.CurrentRenameAction  TTBXItem	TBXItem41Action+NonVisualDataModule.CurrentPropertiesAction  TTBXSeparatorItemTBXSeparatorItem8HintE  TTBXItem	TBXItem30Action%NonVisualDataModule.CurrentCopyAction  TTBXItem	TBXItem31Action&NonVisualDataModule.RemoteCopyToAction  TTBXItem	TBXItem32Action%NonVisualDataModule.CurrentMoveAction  TTBXItem	TBXItem33Action&NonVisualDataModule.RemoteMoveToAction  TTBXItem	TBXItem36ActionNonVisualDataModule.PasteAction  TTBXSeparatorItemTBXSeparatorItem9HintE  TTBXSubmenuItemCustomCommandsMenuAction(NonVisualDataModule.CustomCommandsAction  TTBXSubmenuItemTBXSubmenuItem6Caption&FilnamnHelpKeyword	filenamesHint'Operationer med namn p� vald(a) fil(er) TTBXItem	TBXItem38Action-NonVisualDataModule.FileListToClipboardAction  TTBXItem	TBXItem39Action1NonVisualDataModule.FullFileListToClipboardAction  TTBXItem	TBXItem40Action(NonVisualDataModule.UrlToClipboardAction   TTBXSeparatorItemTBXSeparatorItem1HintE  TTBXItemTBXItem1Action&NonVisualDataModule.CloseSessionAction  TTBXItemTBXItem2Action*NonVisualDataModule.CloseApplicationAction   TTBXSubmenuItemTBXSubmenuItem7Caption
&KommandonHelpKeywordui_explorer_menu#commandsHintAndra kommandon TTBXItem	TBXItem43Action%NonVisualDataModule.SynchronizeAction  TTBXItem	TBXItem44Action)NonVisualDataModule.FullSynchronizeAction  TTBXItemTBXItem3Action#NonVisualDataModule.FindFilesAction  TTBXSubmenuItemQueueSubmenuItemCaption&K�HelpKeywordui_queue#managing_the_queueHintKommandon f�r k�listaOnPopupQueueSubmenuItemPopup TTBXItem	TBXItem46Action#NonVisualDataModule.QueueGoToAction  TTBXSeparatorItemTBXSeparatorItem10HintE  TTBXItem	TBXItem47Action(NonVisualDataModule.QueueItemQueryAction  TTBXItem	TBXItem48Action(NonVisualDataModule.QueueItemErrorAction  TTBXItem	TBXItem49Action)NonVisualDataModule.QueueItemPromptAction  TTBXSeparatorItemTBXSeparatorItem11HintE  TTBXItem	TBXItem50Action*NonVisualDataModule.QueueItemExecuteAction  TTBXItem
TBXItem196Action(NonVisualDataModule.QueueItemPauseAction  TTBXItem
TBXItem197Action)NonVisualDataModule.QueueItemResumeAction  TTBXItem	TBXItem51Action)NonVisualDataModule.QueueItemDeleteAction  TTBXComboBoxItemQueueSpeedComboBoxItemAction(NonVisualDataModule.QueueItemSpeedAction  TTBXSeparatorItemTBXSeparatorItem12HintE  TTBXItem	TBXItem52Action%NonVisualDataModule.QueueItemUpAction  TTBXItem	TBXItem53Action'NonVisualDataModule.QueueItemDownAction  TTBXSeparatorItemTBXSeparatorItem48HintE  TTBXSubmenuItemTBXSubmenuItem13Caption&AllaHelpKeywordui_queue#managing_the_queueHint$Administrationskommandon f�r k�massa TTBXItem
TBXItem198Action'NonVisualDataModule.QueuePauseAllAction  TTBXItem
TBXItem199Action(NonVisualDataModule.QueueResumeAllAction    TTBXSeparatorItemTBXSeparatorItem13HintE  TTBXItemTBXItem5Action+NonVisualDataModule.RemoteAddBookmarkAction  TTBXItemTBXItem6Action/NonVisualDataModule.RemotePathToClipboardAction  TTBXSeparatorItemTBXSeparatorItem2HintE  TTBXItem	TBXItem54Action!NonVisualDataModule.ConsoleAction  TTBXItem	TBXItem55ActionNonVisualDataModule.PuttyAction  TTBXSeparatorItemTBXSeparatorItem14HintE  TTBXItem	TBXItem56Action(NonVisualDataModule.FileSystemInfoAction  TTBXItem	TBXItem57Action%NonVisualDataModule.ClearCachesAction   TTBXSubmenuItemTBXSubmenuItem18Caption&MarkeraHelpKeywordui_explorer_menu#markHintKommandon f�r markera TTBXItem
TBXItem107Action#NonVisualDataModule.SelectOneAction  TTBXItem
TBXItem108Action NonVisualDataModule.SelectAction  TTBXItem
TBXItem109Action"NonVisualDataModule.UnselectAction  TTBXItem
TBXItem110Action#NonVisualDataModule.SelectAllAction  TTBXItem
TBXItem111Action)NonVisualDataModule.InvertSelectionAction  TTBXItem
TBXItem112Action(NonVisualDataModule.ClearSelectionAction  TTBXItem	TBXItem27Action*NonVisualDataModule.RestoreSelectionAction   TTBXSubmenuItemTBXSubmenuItem19CaptionSessionHelpKeywordui_explorer_menu#sessionHintKommandon f�r session TTBXItem
TBXItem113Action$NonVisualDataModule.NewSessionAction  TTBXItem	TBXItem90Action*NonVisualDataModule.DuplicateSessionAction  TTBXSubmenuItemTBXSubmenuItem20Action'NonVisualDataModule.SavedSessionsAction  TTBXSeparatorItemTBXSeparatorItem29HintE  TTBXSubmenuItemTBXSubmenuItem21Action(NonVisualDataModule.OpenedSessionsAction  TTBXItem
TBXItem114Action,NonVisualDataModule.SaveCurrentSessionAction  TTBXItem
TBXItem115Action&NonVisualDataModule.CloseSessionAction   TTBXSubmenuItemTBXSubmenuItem1Caption&VisaHelpKeywordui_explorer_menu#viewHint�ndra layout f�r program TTBXSubmenuItemTBXSubmenuItem2Caption&Verktygsf�ltHelpKeywordui_toolbarsHintVisa/d�lj verktygsf�lt TTBXItemTBXItem7Action-NonVisualDataModule.ExplorerAddressBandAction  TTBXItemTBXItem8Action-NonVisualDataModule.ExplorerToolbarBandAction  TTBXItemTBXItem9Action/NonVisualDataModule.ExplorerSelectionBandAction  TTBXItem	TBXItem10Action-NonVisualDataModule.ExplorerSessionBandAction  TTBXItem	TBXItem11Action1NonVisualDataModule.ExplorerPreferencesBandAction  TTBXItem	TBXItem12Action*NonVisualDataModule.ExplorerSortBandAction  TTBXItem	TBXItem82Action-NonVisualDataModule.ExplorerUpdatesBandAction  TTBXItem	TBXItem83Action.NonVisualDataModule.ExplorerTransferBandAction  TTBXItem	TBXItem28Action4NonVisualDataModule.ExplorerCustomCommandsBandAction  TTBXSeparatorItemTBXSeparatorItem19HintE  TTBXItem	TBXItem92Action&NonVisualDataModule.LockToolbarsAction   TTBXItem	TBXItem13Action#NonVisualDataModule.StatusBarAction  TTBXItem	TBXItem14Action!NonVisualDataModule.ViewLogAction  TTBXSubmenuItemTBXSubmenuItem14Caption&K�HelpKeywordui_queueHintKonfigurera k�lista TTBXItem	TBXItem77Action#NonVisualDataModule.QueueShowAction	RadioItem	  TTBXItem	TBXItem78Action,NonVisualDataModule.QueueHideWhenEmptyAction	RadioItem	  TTBXItem	TBXItem79Action#NonVisualDataModule.QueueHideAction	RadioItem	  TTBXSeparatorItemTBXSeparatorItem21HintE  TTBXItem	TBXItem80Action&NonVisualDataModule.QueueToolbarAction  TTBXSeparatorItemTBXSeparatorItem22HintE  TTBXSubmenuItemTBXSubmenuItem8Action-NonVisualDataModule.QueueCycleOnceEmptyActionDropdownCombo	 TTBXItem
TBXItem222Action,NonVisualDataModule.QueueIdleOnceEmptyAction	RadioItem	  TTBXItem
TBXItem223Action2NonVisualDataModule.QueueDisconnectOnceEmptyAction	RadioItem	  TTBXItem
TBXItem224Action0NonVisualDataModule.QueueShutDownOnceEmptyAction	RadioItem	   TTBXItem	TBXItem81Action*NonVisualDataModule.QueuePreferencesAction   TTBXItem	TBXItem15Action$NonVisualDataModule.RemoteTreeAction  TTBXSeparatorItemTBXSeparatorItem3HintE  TTBXItem	TBXItem16Action%NonVisualDataModule.CurrentIconAction  TTBXItem	TBXItem17Action*NonVisualDataModule.CurrentSmallIconAction  TTBXItem	TBXItem18Action%NonVisualDataModule.CurrentListAction  TTBXItem	TBXItem19Action'NonVisualDataModule.CurrentReportAction  TTBXSeparatorItemTBXSeparatorItem4HintE  TTBXSubmenuItemTBXSubmenuItem15Caption&G� tillHelpKeywordtask_navigateHintG� till katalog TTBXItem	TBXItem84Action'NonVisualDataModule.RemoteOpenDirAction  TTBXSeparatorItemTBXSeparatorItem25HintE  TTBXItem	TBXItem85Action)NonVisualDataModule.RemoteParentDirAction  TTBXItem	TBXItem86Action'NonVisualDataModule.RemoteRootDirAction  TTBXItem	TBXItem87Action'NonVisualDataModule.RemoteHomeDirAction  TTBXSeparatorItemTBXSeparatorItem26HintE  TTBXItem	TBXItem88Action$NonVisualDataModule.RemoteBackAction  TTBXItem	TBXItem89Action'NonVisualDataModule.RemoteForwardAction   TTBXItem	TBXItem20Action'NonVisualDataModule.RemoteRefreshAction  TTBXSubmenuItemTBXSubmenuItem16Caption&SorteraHelpKeywordui_file_panel#sorting_filesHint�ndra filordning i panelen TTBXItem	TBXItem93Action-NonVisualDataModule.RemoteSortAscendingAction  TTBXSeparatorItemTBXSeparatorItem28HintE  TTBXItem	TBXItem94Action*NonVisualDataModule.RemoteSortByNameAction
GroupIndex  TTBXItem	TBXItem95Action)NonVisualDataModule.RemoteSortByExtAction
GroupIndex  TTBXItem
TBXItem132Action*NonVisualDataModule.RemoteSortByTypeAction	RadioItem	  TTBXItem	TBXItem96Action-NonVisualDataModule.RemoteSortByChangedAction
GroupIndex  TTBXItem	TBXItem97Action*NonVisualDataModule.RemoteSortBySizeAction
GroupIndex  TTBXItem	TBXItem98Action,NonVisualDataModule.RemoteSortByRightsAction
GroupIndex  TTBXItem	TBXItem99Action+NonVisualDataModule.RemoteSortByOwnerAction
GroupIndex  TTBXItem
TBXItem100Action+NonVisualDataModule.RemoteSortByGroupAction
GroupIndex   TTBXSubmenuItemTBXSubmenuItem17CaptionVisa &kolumnerHelpKeywordui_file_panel#selecting_columnsHint#V�lj kolumner som ska visas i panel TTBXItem
TBXItem101Action2NonVisualDataModule.ShowHideRemoteNameColumnAction  TTBXItem
TBXItem102Action2NonVisualDataModule.ShowHideRemoteSizeColumnAction  TTBXItem
TBXItem131Action2NonVisualDataModule.ShowHideRemoteTypeColumnAction  TTBXItem
TBXItem103Action5NonVisualDataModule.ShowHideRemoteChangedColumnAction  TTBXItem
TBXItem104Action4NonVisualDataModule.ShowHideRemoteRightsColumnAction  TTBXItem
TBXItem105Action3NonVisualDataModule.ShowHideRemoteOwnerColumnAction  TTBXItem
TBXItem106Action3NonVisualDataModule.ShowHideRemoteGroupColumnAction  TTBXItem	TBXItem76Action8NonVisualDataModule.ShowHideRemoteLinkTargetColumnAction   TTBXItem
TBXItem138Action&NonVisualDataModule.RemoteFilterAction  TTBXSeparatorItemTBXSeparatorItem23HintE  TTBXColorItemColorMenuItemAction#NonVisualDataModule.ColorMenuActionColorclNone TTBXItem
TBXItem216Action&NonVisualDataModule.ColorDefaultAction  TTBXSeparatorItemTBXSeparatorItem50Blank	  TTBXColorPaletteSessionColorPalettePaletteOptionstpoCustomImages OnChangeSessionColorPaletteChange  TTBXSeparatorItemTBXSeparatorItem51HintE  TTBXItem
TBXItem217Action#NonVisualDataModule.ColorPickAction   TTBXSeparatorItemTBXSeparatorItem5HintE  TTBXItem	TBXItem21Action%NonVisualDataModule.PreferencesAction   TTBXSubmenuItemTBXSubmenuItem22Caption&Hj�lpHelpKeywordui_explorer_menu#helpHintHj�lp TTBXItem
TBXItem116Action)NonVisualDataModule.TableOfContentsAction  TTBXSeparatorItemTBXSeparatorItem30HintE  TTBXItem
TBXItem117Action"NonVisualDataModule.HomepageAction  TTBXItem
TBXItem118Action#NonVisualDataModule.ForumPageAction  TTBXItem
TBXItem119Action%NonVisualDataModule.HistoryPageAction  TTBXSeparatorItemTBXSeparatorItem31HintE  TTBXItem
TBXItem120Action)NonVisualDataModule.CheckForUpdatesAction  TTBXSeparatorItemTBXSeparatorItem32HintE  TTBXItem
TBXItem121Action$NonVisualDataModule.DonatePageAction  TTBXSeparatorItemTBXSeparatorItem33HintE  TTBXItem
TBXItem122ActionNonVisualDataModule.AboutAction    TTBXToolbarButtonsToolbarLeft Top1Caption	KommandonDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXSubmenuItem
BackButtonAction$NonVisualDataModule.RemoteBackActionDropdownCombo	  TTBXSubmenuItemForwardButtonAction'NonVisualDataModule.RemoteForwardActionDropdownCombo	  TTBXSeparatorItemTBXSeparatorItem6  TTBXItem	TBXItem23Action)NonVisualDataModule.RemoteParentDirAction  TTBXItem	TBXItem24Action'NonVisualDataModule.RemoteRootDirAction  TTBXItem	TBXItem29Action'NonVisualDataModule.RemoteHomeDirAction  TTBXItem	TBXItem37Action'NonVisualDataModule.RemoteRefreshAction  TTBXSeparatorItemTBXSeparatorItem15  TTBXItem	TBXItem42Action%NonVisualDataModule.CurrentEditAction  TTBXItem	TBXItem45Action%NonVisualDataModule.CurrentOpenAction  TTBXItem	TBXItem58Action'NonVisualDataModule.CurrentDeleteAction  TTBXItem	TBXItem59Action+NonVisualDataModule.CurrentPropertiesAction  TTBXItem	TBXItem60Action'NonVisualDataModule.CurrentRenameAction  TTBXSeparatorItemTBXSeparatorItem16  TTBXItem	TBXItem61Action*NonVisualDataModule.CurrentCreateDirAction  TTBXItem	TBXItem62Action%NonVisualDataModule.AddEditLinkAction  TTBXItem	TBXItem63Action!NonVisualDataModule.ConsoleAction  TTBXItem	TBXItem91ActionNonVisualDataModule.PuttyAction  TTBXSeparatorItemTBXSeparatorItem17  TTBXItem	TBXItem64Action%NonVisualDataModule.SynchronizeAction  TTBXItem	TBXItem65Action)NonVisualDataModule.FullSynchronizeAction  TTBXItem
TBXItem139Action#NonVisualDataModule.FindFilesAction   TTBXToolbarSelectionToolbarLeft TopKCaption	MarkeringDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem	TBXItem66Action NonVisualDataModule.SelectAction  TTBXItem	TBXItem67Action"NonVisualDataModule.UnselectAction  TTBXSeparatorItemTBXSeparatorItem18  TTBXItem	TBXItem68Action#NonVisualDataModule.SelectAllAction  TTBXItem	TBXItem69Action)NonVisualDataModule.InvertSelectionAction  TTBXItem	TBXItem70Action(NonVisualDataModule.ClearSelectionAction  TTBXItem
TBXItem134Action*NonVisualDataModule.RestoreSelectionAction   TTBXToolbarSessionToolbarLeft TopeCaptionSessionDockModedmCannotFloatDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	Stretch	TabOrderOnResizeToolBarResizeOnGetBaseSizeToolbarGetBaseSize TTBXItem
TBXItem123Action$NonVisualDataModule.NewSessionAction  TTBXItem
TBXItem137Action*NonVisualDataModule.DuplicateSessionAction  TTBXSeparatorItemTBXSeparatorItem34  TTBXComboBoxItemSessionCombo	EditWidthrDropDownList	MaxVisibleItems  TTBXItem
TBXItem124Action&NonVisualDataModule.CloseSessionAction  TTBXSeparatorItemTBXSeparatorItem35  TTBXSubmenuItemTBXSubmenuItem23Action'NonVisualDataModule.SavedSessionsActionOptionstboDropdownArrow   TTBXItem
TBXItem125Action,NonVisualDataModule.SaveCurrentSessionAction   TTBXToolbarPreferencesToolbarLeft TopCaptionInst�llningarDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem126Action%NonVisualDataModule.PreferencesAction  TTBXSeparatorItemTBXSeparatorItem36  TTBXSubmenuItemTBXSubmenuItem3Action+NonVisualDataModule.CurrentCycleStyleActionDropdownCombo	 TTBXItem	TBXItem72Action%NonVisualDataModule.CurrentIconAction  TTBXItem	TBXItem73Action*NonVisualDataModule.CurrentSmallIconAction  TTBXItem	TBXItem74Action%NonVisualDataModule.CurrentListAction  TTBXItem	TBXItem75Action'NonVisualDataModule.CurrentReportAction   TTBXItem
TBXItem127Action!NonVisualDataModule.ViewLogAction  TTBXSubmenuItemTBXSubmenuItem24Action)NonVisualDataModule.QueueToggleShowActionDropdownCombo	 TTBXItem
TBXItem128Action#NonVisualDataModule.QueueShowAction	RadioItem	  TTBXItem
TBXItem129Action,NonVisualDataModule.QueueHideWhenEmptyAction	RadioItem	  TTBXItem
TBXItem130Action#NonVisualDataModule.QueueHideAction	RadioItem	   TTBXItem	TBXItem71Action$NonVisualDataModule.RemoteTreeAction   TTBXToolbarSortToolbarLeft Top� CaptionSorteraDockPos DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem145Action.NonVisualDataModule.CurrentSortAscendingAction  TTBXSeparatorItemTBXSeparatorItem40  TTBXItem
TBXItem146Action+NonVisualDataModule.CurrentSortByNameAction  TTBXItem
TBXItem147Action*NonVisualDataModule.CurrentSortByExtAction  TTBXItem
TBXItem133Action*NonVisualDataModule.RemoteSortByTypeAction	RadioItem	  TTBXItem
TBXItem149Action.NonVisualDataModule.CurrentSortByChangedAction  TTBXItem
TBXItem150Action+NonVisualDataModule.CurrentSortBySizeAction  TTBXItem
TBXItem151Action-NonVisualDataModule.CurrentSortByRightsAction  TTBXItem
TBXItem152Action,NonVisualDataModule.CurrentSortByOwnerAction  TTBXItem
TBXItem153Action,NonVisualDataModule.CurrentSortByGroupAction   TTBXToolbarAddressToolbarLeft TopCaptionAdress
DockableTodpTopdpBottom DockModedmCannotFloatDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHint	PopupMenu&NonVisualDataModule.RemoteAddressPopup	ResizableShowHint	Stretch	TabOrderOnResizeToolBarResizeOnGetBaseSizeToolbarGetBaseSize TTBXLabelItemTBXLabelItem1CaptionAdressMargin  TTBXComboBoxItemUnixPathComboBox	EditWidth� OnAcceptTextUnixPathComboBoxAcceptTextOnBeginEditUnixPathComboBoxBeginEdit	ShowImage	MaxVisibleItemsShowListImages	OnAdjustImageIndex"RemotePathComboBoxAdjustImageIndex
OnDrawItemRemotePathComboBoxDrawItemOnItemClickRemotePathComboBoxItemClickOnMeasureWidthRemotePathComboBoxMeasureWidthOnCancelRemotePathComboBoxCancel  TTBXItem	TBXItem22Action'NonVisualDataModule.RemoteOpenDirAction   TTBXToolbarUpdatesToolbarLeft Top� CaptionUppdateringarDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXSubmenuItemTBXSubmenuItem4Action%NonVisualDataModule.ShowUpdatesActionDropdownCombo	 TTBXItem
TBXItem184Action)NonVisualDataModule.CheckForUpdatesAction  TTBXSeparatorItemTBXSeparatorItem46HintE  TTBXItem
TBXItem180Action"NonVisualDataModule.HomepageAction  TTBXItem
TBXItem187Action&NonVisualDataModule.DownloadPageAction  TTBXItem
TBXItem181Action#NonVisualDataModule.ForumPageAction  TTBXItem
TBXItem182Action%NonVisualDataModule.HistoryPageAction  TTBXItem
TBXItem185Action$NonVisualDataModule.DonatePageAction  TTBXSeparatorItemTBXSeparatorItem45HintE  TTBXItem
TBXItem183Action,NonVisualDataModule.UpdatesPreferencesAction    TTBXToolbarTransferToolbarLeft.Top� Caption�verf�ringsinst�llningarDockModedmCannotFloatDockPos,DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	Stretch	TabOrderOnResizeToolBarResizeOnGetBaseSizeToolbarGetBaseSize TTBXDropDownItemTransferDropDown	EditWidthrHint*V�lj f�rinst�llda �verf�ringsinst�llningarDropDownList	 TTBXStringListTransferListMaxVisibleItemsMinWidth^  TTBXLabelItemTransferLabelMarginShowAccelChar  TTBXSeparatorItemTBXSeparatorItem52  TTBXItem
TBXItem189Action,NonVisualDataModule.PresetsPreferencesActionDisplayModenbdmImageAndText    TTBXToolbarCustomCommandsToolbarLeft� Top� CaptionEgna kommandonDockPos� DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder	Visible   �TPanelRemotePanelLeft	Top� WidthnHeight� Constraints.MinHeightdConstraints.MinWidth�  �	TSplitterRemotePanelSplitterHeightdHintPDra f�r att �ndra storlek p� katalogtr�d. Dubbelklicka f�r att d�lja katalogtr�d  �TTBXStatusBarRemoteStatusBarTopmWidthnHeightImagesGlyphsModule.SessionImagesPanelsSizedStretchPriorityTag TextTruncationtwEndEllipsis 	AlignmenttaCenter
ImageIndexMaxSize#Size#Tag  	AlignmenttaCenterMaxSizeFViewPrioritybSizeFTag TextTruncationtwEndEllipsis 	AlignmenttaCenter
ImageIndex MaxSize#Size#Tag  	AlignmenttaCenterMaxSizePViewPrioritycSizePTag TextTruncationtwEndEllipsis  OnPanelDblClickStatusBarPanelDblClick  �TUnixDirViewRemoteDirViewWidth�HeightdOnUpdateStatusBarRemoteDirViewUpdateStatusBarOnPathChangeRemoteDirViewPathChange  �TUnixDriveViewRemoteDriveViewHeightdConstraints.MinWidth(  TTBXDock
BottomDockLeft TopdWidthnHeight	FixAlign	PositiondpBottom   �TPanel
QueuePanelTopSWidth� �	TListView
QueueView2Width�  �TTBXDock	QueueDockWidth�   TTBXDockLeftDockLeft Top� Width	Height� PositiondpLeft  TTBXDock	RightDockLeftwTop� Width	Height� PositiondpRight     TPF0TSelectMaskDialogSelectMaskDialogLeftqTopHelpType	htKeywordHelpKeyword	ui_selectBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSelectXClientHeight� ClientWidthiColor	clBtnFace
ParentFont	OldCreateOrder	OnCloseQueryFormCloseQuery
DesignSizei�  PixelsPerInch`
TextHeight 	TGroupBox	MaskGroupLeftTopWidthYHeight^AnchorsakLeftakTopakRightakBottom TabOrder 
DesignSizeY^  TLabelLabel3LeftTopWidth/HeightCaption	Fil&mask:FocusControlMaskEdit  	TCheckBoxIncludingDirectoriesCheckLeftTop?Width� HeightCaptionInkludera &katalogerTabOrder  THistoryComboBoxMaskEditLeftTop$Width9HeightAutoComplete
ItemHeight	MaxLength�TabOrder Text*.*OnExitMaskEditExit  TStaticTextHintTextLeft� Top@WidthaHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption	Mask&tipsTabOrderTabStop	   TButtonOKBtnLeftmTopmWidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeft� TopmWidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeftTopmWidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrderOnClickHelpButtonClick  TButtonClearButtonLeftTopmWidthKHeightAnchorsakTopakRight Caption&RensaModalResultTabOrderOnClickClearButtonClick      TPF0TSymlinkDialogSymlinkDialogLeft�Top� HelpType	htKeywordHelpKeyword
ui_symlinkBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSymlinkDialogClientHeight� ClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameMS Sans Serif
Font.Style OldCreateOrderPositionpoMainFormCenterOnShowFormShow
DesignSize��  PixelsPerInch`
TextHeight 	TGroupBoxSymlinkGroupLeftTopWidth|Height� AnchorsakLeftakTopakRightakBottom TabOrder 
DesignSize|�   TLabelFileNameLabelLeftTopWidthRHeightCaption&L�nk/genv�g fil:FocusControlFileNameEdit  TLabelLabel1LeftTop@WidtheHeightCaption&Pekar l�nk/genv�g till:FocusControlPointToEdit  TEditFileNameEditLeftTop WidthfHeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder OnChangeControlChange  TEditPointToEditLeftTopPWidthfHeightAnchorsakLeftakTopakRight 	MaxLength� TabOrderOnChangeControlChange  	TCheckBoxSymbolicCheckLeftTopmWidth� HeightCaptionSy&mbolisk l�nkTabOrderOnClickControlChange   TButtonOkButtonLeft� Top� WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top� WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeft8Top� WidthKHeightAnchorsakRightakBottom Caption&Hj�lpTabOrderOnClickHelpButtonClick     TPF0TSynchronizeChecklistDialogSynchronizeChecklistDialogLeft4Top� Width�Height�HelpType	htKeywordHelpKeywordui_synchronize_checklistBorderIconsbiSystemMenu
biMaximizebiHelp CaptionChecklist f�r synkroniseringColor	clBtnFaceConstraints.MinHeight^Constraints.MinWidth|
ParentFont		Icon.Data
~          h     (                                                                                                      �J�W�J�4�b<                           �`-�a�T                                       �l�a                                          �w�Q                                       ��{�R               �f=               �d1�d1����R�>�>�>   ��j�>�g               �,����t�>�>   �>�g�g�g�>               ����m�~[   �>�Z�g�g�d�Z�>               ��a.            �Z�Z�g�R                                    �Z�g�R                                       �d�d�j=                                    �L�g�R                           �c=�xA�]�q�e�U                                                                                                               �  �  �  ��  ��        �  �   �   �  ��  �  �  �  ��  
KeyPreview	OldCreateOrder	PositionpoMainFormCenterOnShowFormShowPixelsPerInch`
TextHeight TPanelPanelLeftKTop WidthtHeight�AlignalRight
BevelOuterbvNoneTabOrder TButtonOkButtonLeftTopWidthdHeightCaptionOKDefault	ModalResultTabOrder   TButtonCancelButtonLeftTop(WidthdHeightCancel	CaptionAvbrytModalResultTabOrder  TButtonCheckAllButtonLeftTop� WidthdHeightCaptionMarkera &allaTabOrderOnClickCheckAllButtonClick  TButtonUncheckAllButtonLeftTop� WidthdHeightCaptionAvmarkera a&llaTabOrderOnClickCheckAllButtonClick  TButtonCheckButtonTagLeftTopvWidthdHeightCaptionMarkeraTabOrderOnClickCheckButtonClick  TButtonUncheckButtonLeftTop� WidthdHeightCaption	AvmarkeraTabOrderOnClickCheckButtonClick  TButton
HelpButtonLeftTopHWidthdHeightCaption&Hj�lpTabOrderOnClickHelpButtonClick  TButtonCustomCommandsButtonTagLeftTopWidthdHeightCaptionEgna ko&mmandonTabOrderOnClickCustomCommandsButtonClick   TIEListViewListViewLeft Top WidthKHeight�AlignalClient
Checkboxes	FullDrag	HideSelectionReadOnly		RowSelect		PopupMenuListViewPopupMenuTabOrder 	ViewStylevsReportOnChangeListViewChange
OnChangingListViewChanging
NortonLikenlOffColumnsCaptionNamn CaptionLokal katalogWidthd 	AlignmenttaRightJustifyCaptionStorlekWidthF Caption�ndradWidthP MaxWidthMinWidthWidth CaptionFj�rrkatalogWidthd 	AlignmenttaRightJustifyCaptionStorlekWidthF Caption�ndradWidthP  OnAdvancedCustomDrawSubItem!ListViewAdvancedCustomDrawSubItem	OnCompareListViewCompareOnContextPopupListViewContextPopupOnSelectItemListViewSelectItemOnSecondaryColumnHeaderListViewSecondaryColumnHeader  
TStatusBar	StatusBarLeft Top�Width�HeightHint5Klicka f�r att markera alla �tg�rder av den h�r typenPanelsStylepsOwnerDrawText$Fullst�ndiga synkroniserings�tg�rderWidth_ StylepsOwnerDrawTextNya lokala filerWidth_ StylepsOwnerDrawTextNya fj�rrfilerWidth_ StylepsOwnerDrawTextUppdaterade lokala filerWidth_ StylepsOwnerDrawTextUppdaterade fj�rrfilerWidth_ StylepsOwnerDrawTextGamla fj�rrfilerWidth_ StylepsOwnerDrawTextGamla lokala filerWidth_ Width2  ParentShowHintShowHint	SimplePanelOnMouseDownStatusBarMouseDownOnMouseMoveStatusBarMouseMoveOnDrawPanelStatusBarDrawPanelOnResizeStatusBarResize  
TImageListActionImagesLefthTophBitmap
&2  IL 	    �������������BM6       6   (   @   0           0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �                                           �                   �                                           �                                                                                                                                             11�   �   �                                                     11�   �   �                                                                                                                                     �   �                                           11� 1��   �   �                               �                 11� 1��   �   �                               �                                                                                             �   �   �                                               11�  c�   �                           �                         11�  c�   �                           �                                                                                             �   �   �   �       �   �   �       �   �                         �   �   �                   �   �                               �   �   �                   �   �                                                                                         �   �3  �3  �3  �3      �3  �3  �3      �3  �3                            �   �   �           �   �                                       �   �   �           �   �                                                                                         �   �3  �3  �3  �3  �3      �3  �3  �3      �3  �3                                �   �   �   �   �                                               �   �   �   �   �                                                                                                 �   �3  �3  �3  �3      �3  �3  �3      �3  �3                                    �   �   �                                                       �   �   �                                                                                                         �   �3  �3  �3      �3  �3  �3      �3  �3                                �   �   �   �   �                                               �   �   �   �   �                                                                                                         �   �3  �3                                                        �   �   �           �   �                                       �   �   �           �   �                                                                                                         �3  �3                                                �   �   �   �                   �   �                           �   �   �   �                   �   �                                                                                                                                                       � 1��   �   �                           �   �                   � 1��   �   �                           �   �                                                                                                                                                 cc�   � cc�                                       �             cc�   � cc�                                       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     MMM MMM MMM MMM MMM MMM MMM MMM MMM MMM                                                                                                                                                                                                                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� MMM                                                                                                                                                                                                                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� MMM                                         3�  3�                                               �   �                                                                      �3  �3                                  ��� ��� ��� ��� MM� ��� ��� ��� ��� ��� ��� MMM                                         3�  3�   �                                       �   �   �                                                                      �3  �3  �                               ��� ��� ��� MM� MM� MM� ��� ��� ��� ��� ��� MMM             3�  3�      3�  3�  3�      3�  3�  3�   �                               �   �   �   �       �   �   �       �   �              �3  �3      �3  �3  �3      �3  �3  �3  �                           ��� ��� MM� MM� ��� MM� MM� ��� ��� ��� ��� MMM             3�  3�      3�  3�  3�      3�  3�  3�  3�   �                       �  3�  3�  3�  3�      3�  3�  3�      3�  3�              �3  �3      �3  �3  �3      �3  �3  �3  �3  �                       ��� ��� ��� ��� ��� ��� MM� ��� ��� ��� ��� MMM             3�  3�      3�  3�  3�      3�  3�  3�  3�  3�   �               �  3�  3�  3�  3�  3�      3�  3�  3�      3�  3�              �3  �3      �3  �3  �3      �3  �3  �3  �3  �3  �                   ��� ��� ��� ��� ��� ��� ��� MM� ��� ��� ��� MMM             3�  3�      3�  3�  3�      3�  3�  3�  3�   �                       �  3�  3�  3�  3�      3�  3�  3�      3�  3�              �3  �3      �3  �3  �3      �3  �3  �3  �3  �                       ��� ��� ��� ��� ��� ��� ��� ��� MM� ��� ��� MMM              �   �       �   �   �       �   �   �   �                               �  3�  3�  3�      3�  3�  3�      3�  3�              �   �       �   �   �       �   �   �   �                           ��� ��� ��� ��� ��� ��� ��� ��� ��� MM� ��� MMM                                          �   �   �                                       �  3�  3�                                                                      �   �   �                               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� MMM                                          �   �                                              3�  3�                                                                      �   �                                   ��� ��� ��� MMM MMM MMM MMM MMM MMM ��� ��� MMM                                                                                                                                                                                                                     ��� ��� MMM ��� ��� ��� ��� MMM ��� ���                                                                                                                                                                                                                                     ��� ��� ��� ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         BM>       >   (   @   0         �                      ���                                                                                                                                 ������  ������  ������  ������  ������  �����  ���  ��?�?  ���  ��?�?  ����  ������  �����  ������  ������  ������  ������������������������?���?��������������������������������?���?���������������?��������������                        
TPopupMenuListViewPopupMenuLefthTopH 	TMenuItem	CheckItemTagCaption&MarkeraOnClickCheckButtonClick  	TMenuItemUncheckItemCaption
&AvmarkeraOnClickCheckButtonClick  	TMenuItemN1Caption-  	TMenuItemSelectAllItemCaption&Markera allaShortCutA@OnClickSelectAllItemClick   TTimerUpdateTimerEnabledIntervaldOnTimerUpdateTimerTimerLefthTop(  
TImageListArrowImagesLeft�TophBitmap
&  IL     �������������BM6       6   (   @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ��� ��� ��� ��� ��� ��� ��� ���                                             ��� ���                                                                                                                                                                             ���                         ���                                         ���         ���                                                                                                                                                                             ���                 ���                                             ���         ���                                                                                                                                                                             ���                 ���                                         ���                 ���                                                                                                                                                                             ���         ���                                             ���                 ���                                                                                                                                                                             ���         ���                                         ���                         ���                                                                                                                                                                             ��� ���                                             ��� ��� ��� ��� ��� ��� ��� ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 BM>       >   (   @            �                       ��� ����    ����    ����    ����    ����    ��    ����    ����    ����    ����    ����    ��    ����    ����    ����    ����                             TPF0TSynchronizeDialogSynchronizeDialogLeftoTop� HelpType	htKeywordHelpKeywordui_keepuptodateBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption"Keep remote directory up to date XClientHeight�ClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameMS Sans Serif
Font.Style 
KeyPreview	OldCreateOrderPositionpoMainFormCenterOnCloseQueryFormCloseQuery	OnKeyDownFormKeyDownOnShowFormShow
DesignSize�� PixelsPerInch`
TextHeight 	TGroupBoxDirectoriesGroupLeftTopWidth}HeightwAnchorsakLeftakTopakRight Caption	KatalogerTabOrder 
DesignSize}w  TLabelLocalDirectoryLabelLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption,Be&vaka f�r�ndringar i den lokala katalogen:FocusControlLocalDirectoryEdit  TLabelRemoteDirectoryLabelLeftTopDWidth
HeightAnchorsakLeftakTopakRight Caption3... och inf�r dessa &automatiskt p� fj�rrkatalogen:FocusControlRemoteDirectoryEdit  THistoryComboBoxRemoteDirectoryEditLeftTopTWidthgHeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeight	MaxLength�TabOrderTextRemoteDirectoryEditOnChangeControlChange  THistoryComboBoxLocalDirectoryEditLeftTop#WidthHeightAutoCompleteAnchorsakLeftakTopakRight 
ItemHeight	MaxLength�TabOrder TextLocalDirectoryEditOnChangeControlChange  TButtonLocalDirectoryBrowseButtonLeft%Top!WidthKHeightAnchorsakTopakRight Caption&Bl�ddra...TabOrderOnClickLocalDirectoryBrowseButtonClick   TButton
StopButtonLeft� Top WidthJHeightCaption&StoppTabOrderOnClickStopButtonClick  TButtonCancelButtonLeft� Top WidthJHeightCancel	CaptionSt�ngModalResultTabOrder  	TGroupBoxOptionsGroupLeftTop� Width}Height_AnchorsakLeftakTopakRight CaptionAlternativ f�r synkroniseringTabOrder
DesignSize}_  	TCheckBoxSynchronizeDeleteCheckLeftTopWidth� HeightCaption&Ta bort filerTabOrder OnClickControlChange  	TCheckBoxSaveSettingsCheckLeftTopDWidth� HeightCaption&Anv�nd &samma inst�llningar n�sta g�ngTabOrderOnClickControlChange  	TCheckBoxSynchronizeExistingOnlyCheckLeft� TopWidth� HeightAnchorsakLeftakTopakRight CaptionBara &existerande filerTabOrderOnClickControlChange  	TCheckBoxSynchronizeRecursiveCheckLeftTop,Width� HeightCaption&Uppdatera underkatalogerTabOrderOnClickControlChange  TGrayedCheckBoxSynchronizeSynchronizeCheckLeft� TopDWidth� HeightAllowGrayed	AnchorsakLeftakTopakRight CaptionSynkronisera vid s&tartTabOrderOnClickControlChange  	TCheckBoxSynchronizeSelectedOnlyCheckLeft� Top,Width� HeightCaption&Bara markerade filerTabOrderOnClickControlChange   TButtonStartButtonLeft� Top WidthJHeightAnchorsakTopakRight Caption&StartDefault	TabOrderOnClickStartButtonClick  TButtonMinimizeButtonLeft� Top WidthJHeightAnchorsakTopakRight Caption	&MinimeraTabOrderOnClickMinimizeButtonClick  TButtonTransferSettingsButtonLeftTop Width� HeightCaption�ver&f�ringsinst�llningarTabOrderOnClickTransferSettingsButtonClick  	TGroupBoxCopyParamGroupLeftTop� Width}Height2Caption�verf�ringsinst�llningarTabOrderOnContextPopupCopyParamGroupContextPopup
OnDblClickCopyParamGroupDblClick
DesignSize}2  TLabelCopyParamLabelLeftTopWidthoHeightAnchorsakLeftakTopakRightakBottom AutoSizeCaptionCopyParamLabelWordWrap	
OnDblClickCopyParamGroupDblClick   TButton
HelpButtonLeft9Top WidthKHeightAnchorsakTopakRight Caption&Hj�lpTabOrderOnClickHelpButtonClick  TPanelLogPanelLeft TopAWidth�HeightdAlignalBottom
BevelOuterbvNoneTabOrder	
DesignSize�d  	TListViewLogViewLeftTopWidth|HeightZAnchorsakLeftakTopakRightakBottom ColumnsWidth�	WidthType�  Width�	WidthType�   
Items.Data
:   :          ��������       20:30:45 PMDetected change��ReadOnly		RowSelect	ShowColumnHeadersTabOrder 	ViewStylevsReport	OnKeyDownLogViewKeyDown     TPF0TSynchronizeProgressFormSynchronizeProgressFormLeftOTopBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSynchronization XClientHeightClientWidthrColor	clBtnFace
ParentFont	OldCreateOrderPositionpoMainFormCenter
DesignSizer PixelsPerInch`
TextHeight TLabelLabel1LeftTop	WidthHeightCaptionLokal:  TLabelLabel2LeftTopWidth(HeightCaptionFj�rr:  
TPathLabelRemoteDirectoryLabelLeftXTopWidthHeightUnixPath	IndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  
TPathLabelLocalDirectoryLabelLeftXTop	WidthHeightIndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TLabelStartTimeLabelLeftXTop1WidthQHeightAutoSizeCaption00:00:00  TLabelLabel4LeftTop1Width/HeightCaptionStartad:  TLabelLabel3LeftTopEWidthBHeightCaptionF�rfluten tid:  TLabelTimeElapsedLabelLeftXTopEWidthOHeightAutoSizeCaption00:00:00  TButtonCancelButtonLeftiTop]WidthIHeightAnchorsakLeftakBottom CaptionAvbrytTabOrder OnClickCancelButtonClick  TButtonMinimizeButtonLeft� Top]WidthIHeightAnchorsakTopakRight Caption	&MinimeraTabOrderOnClickMinimizeButtonClick  TTimerUpdateTimerEnabledOnTimerUpdateTimerTimerLeft)TopY           @   4        �      D4   V S _ V E R S I O N _ I N F O     ���   6                                     �    S t r i n g F i l e I n f o   ~    0 4 1 D 0 4 e 4   >   C o m p a n y N a m e     M a r t i n   P r i k r y l     n #  F i l e D e s c r i p t i o n     S w e d i s h   t r a n s l a t i o n   o f   W i n S C P   ( S V )     *   F i l e V e r s i o n     1 . 5 4     � 3  L e g a l C o p y r i g h t   ( c )   2 0 0 3 - 2 0 0 9   A n d r e a s   P e t t e r s s o n   a n d   R e n �   F i c h t e r     < 
  O r i g i n a l F i l e n a m e   W i n S C P . s v   4   P r o d u c t V e r s i o n   4 . 3 . 2 . 0   6   W W W     h t t p : / / w i n s c p . n e t /     (   L a n g N a m e   S w e d i s h   .   P r o d u c t N a m e     W i n S C P     D     V a r F i l e I n f o     $    T r a n s l a t i o n     �                                                                                                                                                                                                                                    